`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
o/j/gktqITv342k9c4N6gVY5MXOc6DIxRLniin5L9G2M2MclC78EfGauRJw+XLAsBJXuxpH2WKpY
oKng13cMVg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJBnQK71+BNUyPq0WjI2RfQgBpA9+MXxZklWXl3WPdstyjmbVaqIwTQl1+lYHmf6dhiSx+cInE3d
+P6kTNovtVAa3ICJzhd+egPNsUXfKFzR394ry9JasOskjMjk7yekZuA00KONTIjMGQdm4ar8u1Py
XirlobPNM6/c5Cv6LKw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Igb0qMFSkLXDt+WWNCwf+iXXyT3wugsR+f40LmORXEVd2datRoJkU9PgZnwNYJv6bvSwNdB3edLI
YHH4hq0BzgdhvEzfPD14btMhdjGbj9M4ExXVWDGjW2P+QutLmLcZMkKvoAsr/E5K7SPPMdFaqn4+
ez0NKiAhWRlc1TmQc9TbL0ZsBkOtRw6gDYruhxEQmMYGOSjGh4b8aMLmZcRUSds/FzsMfHMkXRW3
ZLSubU7ai6+X5Putvd7vrhBeahRThV6I0Lf2JRFIbZu5rUUs5ai2IrFSgIFQdIvMB5rKRI5QjLyr
k4BkJWvJujBOLXyY/x+pGnDc4V8yJD6wXdSnVA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I5VzaK2qu2FJmXT3xhqIDN/KQSXsrW3nb9S0LhCJP/fMe/1Ojthkn3n9b2wgOQBrYXLiP/t+ZS6c
Q/fAgWmkp68jcBASHbsycHnPX5j93TAYDvH6R5NqmRzcU05DKjdKkqtHol39+NaEeX1f8nDC/F1B
6zf7robWLOTAH9K3akfp/4TpAS+scwidmr/o547nsuQYB+45HsEmIQJyxACFKjJxY6ahbKyDC22S
v6C68SiOef7eu4rWrW462RYSLpwwOQKo5vbBhhXREMHyCMcg11eveeeSlOwQFy/mSyxBTcCcYLRm
YkGk0LZU281pxtgk4S4hkVQLT0p5sMsjoIrCLg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HSMYftaO0K2A7/2vhvca0OnylUzUn+mNRr1j3Ee7E+AF4UbrbDV2Cw0oasQVKVKNdUByWnWF3aHP
0ts3kvG3f8Snqe2cAFFWXam3erR2Rj6xrytp/JfvNXIBQFOKpQAMZCC6bM2CFoszG64k+uJTc0by
2fDE0UHTSuz9chEnJ9Vy6LcKH0qI0p9IcYN1ePOHKGjQqhJM0BN8fJo69vwSkSxoAdyB5o7va14v
7tR7eE34OtTwDXZCMZk5f+Phd75JALwmuVXncU7M5S2WnyPslU3sVJcnch7aF4sljZVhI1FpoWKt
KVhgK4spijPbvjXcDSkc7dCDUh/Wj04GpE+vLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d0aYonu/bykDRb7euHIzCz5mWCNmaSle6Mbq0GKaQNyJfjs0qavqNm1V7xFEGDIdkZC7rR24uRxK
b1k6uDweBU2VM8fF/sJtf0w2MOmILLA80RIm/uluHdREzyEaGkx0rsnv8MbjUUecWLWvGfitpg4N
Sl8r6y5KIa4rzSAoOOA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lCKmNYKFTYrMxzL7QW9Sg63joGS1FWrVke09b7jmQskn+j2WW2yrlJHWc2G60QvNwxv6fWPvwVkE
t4xod74PA6h27LPvWuXcOc9YJue+DobGI96k7chBfpY4A2IY380BpaNUY2lgsgrBi93c+YHKs7cT
j7+aSZMLKZupjghs/572g5jC0gXIyW8PxwMptlBHhakXttaIAhIcNopify6N7jag+h1vOypGANJC
DeMz2RK50tD8YG2LLTVlzDU2t/r0EU14fFTRxZDaLMWy8SV+4pXoISsgIDm4wM74Gx9CwIrv3kpE
OsFlJ8QsM6CrCRyX40sji7N0pzzX4k7akuGShQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 610096)
`protect data_block
fqX53hEyvx0OcSsEOHxTipYLDykiOQuiXtpFhQFKD+lgKj+lNmwxKzm0nXcon5KurqnuWx31B1AP
ZezKdSuFn82bA81YDiGfH5mD89eq4B2pGvfKYI5bhdh2Med8eT2fc5VSyqz8TrIDbtH5Nt1NsMki
qqnSfUCyhyGqDMG+nLItCB7fi6qgz3uaj5G4pRhYTsKrtj0Jmew3JI59Dni2d5mtIMeL+FhQXre0
Ef0LJmed1HlRpLQPzGQ5hGTAstCor7daZ2wMFSYyysTvapmsKgym/TghKx0Haf7a2+TdGaDF5iMw
Us0ZTt2Hby4Hixk8+4Lmf6uh3E8ck7SxijqObRT/lh6TjZ4GtZTG5WGb/feXRAI8jgUOhGzS0+Ul
nf2tBkpQb1AO4s7j05PBmbIT0y0vW1g1CGwuALHFVqgDdAQvClnXgNcXqS7l+D4ThSoWIiy4Dpws
xy8pXaygBkGQRC21uFsNGtO85vQfngAPsAzU7CALdQVU4n/5C9uVexLnXsk+C/9PYfzkgQtfipWb
N5HfKRsIims8nRN0t3hp6CqX8qpSx6FXd8gQNYvyTN3W5b+xPm7M2/hY+wab3kWwnrcQfiQgvbWe
v310MHHwk9MeuL2C69NnmQPzsc0Y5Jf98kn4b9oAKztifSA7xeemxpIsBN2o86g5l3v6W9hIBoa2
NaoAURgVsc4ZlvHW0h4GNTwjPJeOteCfD4ViPFHi6kFXoHbQGwq0M9999hXbjomSIYNuCEulLpHH
mOfSntj9Qrqdw3DrAHEjuVHSsIWuDM1+d0pxbxmc2B6Zric+PtrPT5PxWLUF+iG7duFeons56vcQ
Z0n4FztHdaud3lGFCU8Ql4k8Z1kLew31ebG4bklQprekXkgoKFIey9IpyJr0Wziqn/nqfzeh1hl9
s4gANEHjLJfNLHdzvmffEWY1LSCG+r85vFnbeKul+SJFGSSzciO17YF07L/Zo9Zg60mjVbB+n7KR
daAFwqvzSAmG7wyUohsEXxZa31l4Rd4tXijzFnKznv91GA1HhauAJkTlU5SQRFAS36qm0BiU4JAM
6QWKF08i4ABxRo8g5lvPrJ57GTNsRf58aw4ogBanU5b7nxzmp1ajalKw7nAoZiJuWcFjm3o5S2Ak
WQkyVAGIwmcfuHAIWU/kdRvmcnbu35YsCP5WIY32aniKeK7u8lm4K3HuBjUKqtJB1pBJ257g5swf
p6KU9XfAFOTGRRRV976JmLLFvzVADlJihqgT3tWrfkTn/vmtjeL6U/PWmxHKomn2MLZ74DKw6svx
hILbyCdHhji277M/vwRAMVXc+IYR+Bnq+KVwW+Qtnf9Nw61Kt0x+iP5JygLUGm/p9md8P4OmjAIg
tmhfkKgBZJvlI5dH4NViWozC4KlU2gNneV0XK8Ns+HY+OuD9kyWc6rlkOc7BDdY1tRrJpjYAIhIY
CamxmzgkAP/fLrfbC0hI6WvvistE7j4upJu+Gn3Ts2XslgAHXu9Ih/BuxTL5DDDD65/dcEKo3Jij
mQ5YdElWFyHWK2p7Gs4nmIb0nBf/qWO2/01FMBubg1ZC0Td27SI7SiITDWHUvilnKkGkk6gDT56P
sjCtSISuj+C7aTCO5XesEOoahs3xEg1V0AttsPWSDiMBGVLBke5PJPtxUi8RSFPDh1LpW0WG8Qz2
XXe1vq+d/pd6vmwDY8f8Pygj99UBmW+aJ+X3Rz6fQjY2iDeJBI6zramV1qEyKKRpmeMlo0k7g+H9
XlXVer1aGYy06PY+aptTlspJ8vF/32ZOvEDmzOrsnqW1Vaa7GCP6DSEtn7wkNc0s4yOuFsCI+5vf
VCqkWA6Ot2w79zUc75fiKU82LV6WFxXnFLJhQ3E4AfdwUYgzGXbXy6kjEaLEzJJy3uqoEnUuzp2s
//g+9BglmSb3CZHbpqcY7aIwY1tToJHsQ4M0Sj8xeOBlw8f9eRwKZJZGj419qeEvtQ3y5HBLLyi/
MGCh6n27TJiagbbfjy/XspNq2R0kHTmoGB/wXJfEFDichC3QS6/5Q5wrOvpK8h9FuT1NBnDCBrU0
qjsO9WcovFXj8qKNc3xiPsC9llNHN7o7g1FN5H3GVt+cUHKH3iUYWMu/J91KBJHbi/NuhEbWbRBu
KAz2MOVQ/v3BYTDgSy5Gx4wGLlZYqnsG8bC6bcYiBKsFceek0dsEb6IlmU2m1bXoEr0cAUta0UGm
Qh/q3Givu9dDW2lwYE+wekUPLT3rARsEMgh/XGUqRrktg+xeOW8S9gEoKU0Qzp4FBNEMb/rHcyz6
1ZC7zecLxKsXotwJwF87nnwEeE6wyidULvAekcwVkNpeonB7EjrpWNy1f7ZO6XC36rePkXyD7qg2
fHaHNCs0bh5wthUO+CCpByZ9UkJwwsTIqr+dPguiOQ731jieNK/WjiZ74onmZjK4eRQxwPFdt6Vp
4HHBm42yfyZwfdnf89m3rJJwWfTNz8Yu/ROMHuNcqVAxl5sJiBilML0QO3mxdqUwNGUpNEZdPXgp
y/2MiwJ8QV1nifpUoK0Njyga+H8fndUoSJzlp1QBhh9/yHpSScqCpD8r/lyJIgkdBgoRgkYe2n4z
Xe+vuXq5vQ5Dt0Pf/8qwi1SNTo7wwwK6u/XRHPegHZKafmHijoTNDkfIafAM66CGx60q5mSSMRGv
5MIwr+vatQ59HIXBrezGhGU/+4jL88AGvwf25b+TjX7lkwL1lN+A1se57Jbkmo4gd0ZEQtJ9ke1M
BkK3wWiRtFvcw+1ithkrNSwYlTDtwpRbqmn4S5SutvotErUd9PX39FuZ/k2rhW6vkWxJF0J80I6J
iWdqtmK7miH11/O+2NGGiE+3vCS+RJKeRWXRXPGP2jtTqZtUEUT8fQfCmdKg3bN6VOIVcbXIugIu
7JBEK0B0ELCurSo76UlA2ZxZekjkL6I20Zld8SJhlGY4OM2Rg6N5FG6ofpbL578L/TS+DvEkJxDK
TzxmXr+m1Ew2o25DkEjua1WtzoFaX3TLehgMY0pZsU5hIiGhlbF9oxQ4CsLx5lH3IAljNgZ+J0aZ
fKduO1VZZizCZeU74YN19kfMG9QmPkUY03KVRMSxr1Aavlj6HR2I+sa45PYW/CEmdIFoipZug9Lh
L94Pp8m7ggQhW4aQIhf+BFoZ5CXpZ/X/vKuA0tiU+NhIJop92sMU8JrPJYc+/KZnGj2Atvoo4Z+E
QDE+ANsfnGlmMK5tjH8IBTMvzqYQZP1Pisipo5W6icoZu3tTS+VjXnc7JrBNdLXtxle2Jdev7Fy2
hMmXCpmjEyvES1UfFm1WvpbbS0tfpL40PXEPMztkWKYXcNBLztVgn4xYJkjd0PIuw3RCJFh9a58+
gM2eVEwaXwOcOrb1JY7ahMIFl8Tz2Gz0uajXsKpHRY2wALUxsFExSECNX5K8zfOo6Ie2/5Avkgg8
o0k5R8KyKRhxzUT4KIlm3/q4/60tGhxLoNIAmu9uJdqzLABAHhjPzIwuQKtB10Yt473AU/M7BUYj
Oc+uN8UVzf2tncLD1CeOOcpGpX6M/FKS3j+mmMAkReBnCnLnAzcHTjIATHV6Ljeore/ctjplYWBL
FHhwBoYtk5zuVcHqF/oVrr0ZPmZ/YWBTunvf7ughiU/dOi4Mls2epbtrysf3uTa+PVSys4T9hx4c
K4kc2S0kEI53x7HHcW23NTLwikBjUP7/nwglzg8OtlgPMsppueXwrQJczVr0ziPsEUzf0SqainoQ
W84yUvvGATPKUZJDTUTNCx5EASwqn6uQ4I9wBP8CcC6YsQBFDdRR3vXwMEogocwVwLW9R7ccLof3
nKxZvHv23s10ytPirzJenBWWc2fkR0iOF8gN2nxPWVrE+OpbGrym0t1q3VFlGN2+YmNICejmfblL
eF4XlXcoF0n6hAoScANgNjVbbUcbO5URCT5bk+dJ6Uxlp63ILaiWUsNVFPsKbNYTkQw3DUPYiWv8
0r0NlO8mUlyMOhjmpf8+dS7FeGVxPAuTAAmUq+xYVy95Kzov8hME8k4ajuXp/8609NdunDq6G/fp
/tPKZ0ehTkELYELD8ghRs/7YFq3oFFAIUFPlWqJoiNIJBmXEckw7lFxFVsQsb9l5X0VZal15sxPh
hnEwLcNO3Fk4wt2nBMezuI5ggxu4tyrWIbpE4tHdMrQopw0da71peBJXhCtGTw3dYS5dS6SH911s
y4Rc5IHFZj5jMbHwtb1N9Hq/xHKxdBF0kFymU6o0MOdN6X0ZVqnIwif7bvkZR0FuhcxEwhXVZadu
LM7Ht6rT27uul45EwYxSxG1TKeQCpi9+4X/IiIKa+eDV4kOPPPsjOmEzcN4MnrRA/MtX96BKLbw1
Tgo5FS7FzGayXFeF6j0hykw59e06OizjffDZd6nMmJjOWkeTMiHwnuPTflp0Lb1N+NlN6gLCCSjh
4umBt/gQiI6qKXT2mki4J3isBHvaB9Iw0JYycBvRMyetHvh3/YU8XKOEY6dRUca2JXr3OCfrm4rn
zvpHsFPJ2mPqmbWnjaz3uT2vkVckhMi450/1Q+NUhAHT467TavISRYhMJjIAFKKGTlf98t4m7E9o
zPYZdPRyDjR/6rpSUINjxWXyYGZTtNmeO+chQSWVv3jTFCzIdy8Z97KJWWqjsJ/X3M9Yw/BWN4w6
rlTnHzAmFwiYzrjz89DcN9dov1QJtgh0FlSynUtD7Tzk7+kuw3Kf4JMBtOeRnAiWrZJQci0TAylY
wZHN9j1lTGe94cE5sRpC9d8fOtOBsUDDupNtxYsiany93iGz8BS75wSvLUwG9U2+0b/BpppcVyYK
HQ1YSELh14FUAxfILcp0DArFSPmM3fPpAeXFyIyvN2KK6QkQ70OFZbfQefivuOI1Wj1kYnJSkCE+
9qLbrEh7UaMYHmOBl9u1UJe29PBMzTVaupT7cx9S/locRndydGLF1q1v23EPvoy/XWmu1xB71ITU
XQQqiAEgCsOsCSiBfYj5wrwSzcGyxiP6qC3FVW6IuUhJSVjtUPwyungXZfQeXJYFAnnC5o8efAnj
2jFvpFqLX66COhCbOj2U+DuatBRIrxKPRqX5ro4SX7nYZY2TEs4p5UpWQRTBGyPWspSGjDWr4THj
0HW/bc3eKvL8wybRFoKI6qLbMmh3K4C9pZL3icidMPBe3ipUc7d1E25Mp4F5pLnLYZ7n342R1DUv
LKPjdDdRxdZuJk8GUrhLfn5CCylpHzstd70vSpjFpV913DkFMp9fSCU8rRjtbP4O7o9YRx8+XdNe
PC117Ncx+UpU6UNwaKuQqMMF3wQPcJn4C2VX7fw0wgrzzi4xfeUVAwDxgfvub9fqDBMJn8Ypkl39
lrPUzf3flETqIgs7N1x/CV//Wvvb4yJtlo2NV1qhyX9gq33sUMnjvWOUlwI6YFhOF64TRoEoHt0C
PsiM7+RQhyRQe8ZiVsyBlpPlPf/GarSMb8gVtiseZ5ftgI1oAwlSwuJRUgHFCP/rLWjKTqji9C++
DLzo2coJmCr6GSpkxL4UTrzWFbKrg/QcUrbW4+p1ivixKa+Ao+OiVHgYDb8APxBsYGqFCi2Kj5wf
aJo0lfGc1fkKDPpaweiza5Mri9o0kcLnbbeG605Lzl1NMZlx6DFiQbMnALYB0q2NOyzdLPN/eUDv
20DTJoKJYDGSpVYs9m8yoFmA9SxICCNWFWbimejnk7JdYyjaklpOP52cW3/4xNk1UmESUME/3ohC
lB+qj94YaeoYDt1oCC+BaHyWahwcWZr3C6w8AD1huKoMzqrBJTeDxbhBMJa+v6+YGuYQVHztNwVX
mb61t/pd6qKmGl+Ye8DtqO477b8b5V5iqQtpgA+IESrJNufQ1XV5l3JIBmV/tRPHKU7th41kFkdW
HfAUZxjby6B+4MfzwHI1GxE1+v5Sg457PGlGKRWJALStAmQ2ya1LIBRQj1dyzRML6Wn7sxhg7Ebo
v1N572pRcsKe2h2JHzMZ1zMWeziSKtmtnkNKgfcnjg1bPWm/rwuM1t5o+isu6R9Jf4/qK9GS51Ko
M7ExscLAW/1kZJX7JrXTeeLye43eWJTS9Sm18QCxXWfLKkN5Bk/LW7pFS/mDzUpOhFVSNFkD+BpG
MWBhWjbgXWjsqj7D3jD/K+MhCJh2XhmZYGhdeoNxWjNAwG09etk3ciIzEdzJdV9pps+xiYMY4Quf
NO+HAc1hntKF2hiiUFqJu9MsQJk6A7ZFOTwF1PzVjnKHIPP/omBZHqtcTnjqoy7ajnrOuLwzZZOK
eZ+nR5PIUNHnmtHkkVafOyEYEsuVBIPN6I1xfilQwqnW+PrWtjnYN2EJvvdihQwKhN4WyLtdvZYn
rsx6WVs54CJhcxZaBvH7wcvkHYBSMmz98sUWoTRNLcA63q3oAqTquzmhQF7bGrrXHLywrD9wutj7
l9lzTgSxb9pKeV9PSt5bOe62Xkv4XSXbxxnIQwMxI7mtTbBtsXp293TwPnERajZTFMjnzgPfrHI/
D0f0RzgQ9tl6IssOfrZk5hzzJiJ8BNUQE6++WDRbL9yqtOm9Bdj+5nU4QQnmI8C9niarGVXfMUVu
2oZjTDT9F4iP3AkyCkQjoMygkMYKj04sAOge3QBeKY0XM6dLvVAU0eaBimMfDKeHT0gV34wio430
mfzaR5rgYr78LT+wYXo6YbTdjgl/j9iqb1N8AeRKsLW4Ovsda4wOmCSsPZRbIgP+fODJSqim5P8U
ausSYLJYexvSIdX33k5fcW/Dty2OO4H8qnGrgOYQQsFu/AC7eQozHGy2SDqNvS/t0JKS1aBRnySJ
4te+ZUlFe7BqCXictt1N2Ark8wOZNSh2RPoTZdWGzZyQrkKpcqF1aUtgRwYx6p+Ihb0C0Zt2h7kF
cqQQYg5EYhV3KTxVar8loohBtep6Y4N8OQkZ2ocatWsXxN3llcttEsR+vp3ioxbWkV7iEc9yeDMi
ES0mZlrO7NMdHBIXU6tDD+xGVIA940qPuf5gPRVoFJsVc/d8jj0MDs8DhWXev+UsFGrZOaKIL780
HU6Ntt8jIIBP/4BvqkVLCJgXUaCMcRhZ/lScMolXdx3YUzKFnA26cO/q22crL0SWmcOMQ45a2fN2
Dq2iA8eEGl1lsbgXmVIm6uWib0PDLAqKVDBup5EYfwOjHb+tyBgu4O4kBTaUKFdR42PUQwl+GT4F
s1lDpEAbtBJzrdk9HJBs1E89qlnqxSfTpCwzqSAyCgNwgFlYj1mtGfJ/qsFqMPn1gZJEP2ALKSiu
Qyc2JHBB6WPIm0jtsZf6zrotKPcG0rv/HhVxsiiSC7tN2P7pI7KACbegc7xHKomuemXRcpt6XeU1
DNv3xCfCw7iFr6Aj8SUDsT9dU+f6b4UvZc6EHt6yiAI+2DjZ8eHZ0+bMgxEv2WSko0E4tWiuz9V8
tEGHNygnH7XVVou+UWWZo5nSwmokieWo7u0cRt7XGfz6t06oWZlV6kJPzM/fwYpAG5sgVVg+OoPl
pVQwoJb/VfDhjYm+uosFwLtP1XsH7S9VUZrnhgF6KaN6ovGb3tIsw6AQ1uO0ogHylDsLLyTDEwpN
TH/n7Zh/7ynvorNgPUqAxvnqEVM7c29AhVOEZSaUe9ATGEVbv2jMSQL4a53/EDzbhFc1QwB4FDDB
llwEIPiZ3sHrmbW//tlJxzE/psSFBHzbeEMyOaq61GM1su2ul6O0Kj9sXMtjRs2YwLy8ZnId7yg1
Wks9vzJH1sJLNZ61GZfZbj6vXp18sLQZw+VUnuh1a86U4H7tAzoxZc9BZuCZrmXIE7caeU71CXDX
EafrVB+L0F0triHueM0K8q3Z82GlTLTEiGfRiVzVRGesAtNWhfd+m5IRP6X9HHV3QpAoh/Boxpb4
PPkpMoQHK9JbxoJ9kKvUWfjDotyoz/q8hd0M579CyvwkwOB8cyLFbPuxZmCv+bQrAJET/5y1Lldc
XY7aluK2OSdN+2TH9KXr7PrCYY0j6P9QXEvqT7l5xg3JFzpRRKr5EZt5oYMpk1vtcI/0GeTtao1R
sp/Mtxs58zakWowSMYCsfl0oACkd3ahSlyo1Yes3ke69HRhKjnIeNb5tCXSmfA0FLJc1x3exOeiq
sMD1LnMvYOg33Qxq5yLCgRfBU5oVkiCy8+A//r+LD0vGm/EaY7DM2RsMEy+uxZV2mDFa1BuYHIRs
wHY5BdyXT2zUfw7JlZkBCYDs5KYeR8U6eWCR45erfHZPREBHwsN4i5+tRp8XOjFNVBgVmq/Ad6Ne
4NOCXRwQ8pBjmsP7kyruEo8XDa60rJTwp8SIKgd78Ky01qRpNn/qautVlIht6OC92mW0TtDZ8t/j
sEmpCJDsv9EkzpArXANtcesRrgaGThDNmDANuNJcENCH0YklshsFNFGovXQQC54K6pKZMnLjm8ua
D7z+P4hvkGC+yltCABaqf45TlshuWBbLo1lWwLvfHM1WuJtxvcUcSsaGNifxO7tmLgBUMzLqHMJG
5vp2kfBHOPOTMugk+E1BykzYmJwQSTli9lbuePN0abb+QJTBVx+5KTLzHMIbGdKEjzezWlqsyyCF
BNFxz+cd2ckUmZZaAsc5/tMgMT1gSXtrttH3ANGkVohz40ilcCPjxSxPe0ECPmtLk7om2hbz5aES
dG22GQyMjjKQNu5SdDIfqYVTt4oM+7E2epV/TzyCUV2sJlKvMJaZkRZVInGmSMzK0zvju4QyrLiX
w8W8WzbdpXIbG0VGpMUi5BFe+XWOHqul/R9LLVG26Fx8foQruUcooSIADDibfS8lPDyDfwQK2dpM
8XcdMRnkBmVuI96dpN2/15E2PtzegB8Aihz/R90bin+MzUnfdCJxpJkbTrMS0siuwZOLqETfbg91
y1TgBSK74I+CgsaxohaiTdDhrtD+WYmBUqlh1/+5E4UMMQTbM31ayRYMZUlK3zec8KFNU33JuQ8d
xJD+FYjskbH//Am4pzRV3voNI+oQXSlxZN1sLqLo2sB4pAC30S5eeX3bsUuap++HMPLB3TAqsM9c
pSq9LAFWx5UgavHTBHFm5w7SU+H6xLb2S8FY65+Pl5zWUcrKMAs+GwMpKYkpe3xSJnSl9+LSRwJG
AwkWBWbKfMhOD2DsNJLcBP9xXhsUpC70swBcJx6SNNanOWQ3n+WXcKcSh+FwaMU1lebxTdJOgP+Z
7PU88gtyD+++wYv7BPC+sToyk2KtI6PjSnUSnVtXLsx8iTh/Jt6gn/olbaYibTyx7Jbl3miyOEct
vUu0yD1EYetgq0BW+M6QHq1OWpCSuNpNsblSyJfSOxVZ1ms9l1uYpnSWMbx0lVfB1crfYSkT0Rub
owegqWH2p1QdifdCteLncTcv1OEY8G0bL7qSHACNnWq5hoGk70z+CPLU06bJGGhSqOCoKfCssBg/
k/yYCtqbbgXSoAGbgnjm/OCJWialv6izW9SHekRe8jf1TIEqpj3wZ/38obWatYIuDjhlQhBnsUOL
gD6YaYY9krw09jCXVDvnTXtpCpRgJ+CPeL7gyZocoEqHEVJSuUohyR0P6mhgcDjbOshO9NwMDoRt
7foRAiNeLWCoDnsox3HZtCTUQPSXsJqvXWcQQbKCt+3rSuiirucaRGARPx9zB15RR/JM6M0+iDHs
2toIpCZccw8LWB6BJugZwFkismuGunGMVa+W9P2d/0uY5NE9r9kwzkeFRjVciqOwhyStYOQpiUpl
gFwcNcp6wQDwPx5TtxdO3fiEIIYkcSIz11gXs3e2hkt2CDQWsGRQ5f9PNOmPLymgsTtoc+rqnDis
DzRKvzMIJcBHvT7yDl7sZ/DvdHgju7edcLO9DaCFAb6PztPtg43P0RciE2L8uLf9Tm5p4Teviatc
0NsirWlWiKg3JDMIrQYEjozO8SV5SqVdBLqMsVLE4WRTdLCbvC/myMq0htcwOm18EQLo8G/Jke7N
i1XjPTBohRT3vFZteRXVCmGtYDjQNyfAS6u5eTiDTnQkFNpuVG8LeXQ0A8Es7QzY9sqGHZJU4FZc
qadxgElB3F7uzAMkLg2L4CKK3Qi/8rzP0TUEr2vp66lvWh1Kf/87P5IsNCdCXbhQzrRbPiVVnAWL
dG9p+pZSawUpjMB6TQ0z0a++hKo+G4tVPIAB3lvF2TOycEnCyDFTQQ1dtr4XOMP37zrDPF8f54jW
jYdN+5Q9FZRmEhMYMXmnu2on9DfUuWv+kcPmfoaVpND44sWfOlpP6WdoKhtQeYAU9+1hyLYx7LDM
4NQHKBV3Nn9zRJM+Hqv+uvDmE82HLwmG+bgTPxnIa97zKkcKrz7rWf6XpRtiE/58NqSyp4J3waRc
2j8i3N2KZUyhT2mMGWwB/1IeKyG8wpIqRN+sb3RebIzVLBWjqTAti9wxOJEbsXHA3cRPgC7v4+xH
PLcIM9imZEbN4A422wgjFNc2lR3MmZOIMSFNnrSDsaoS9U4hrRKc4ZaR/+ev/1fTSkgcSk0l73I9
Gu3FHlsLLTo+W0Qewok0qpQnRCm08FIhOVCgzqqUv4CYglGKydRlYMT2yE7kNVjH23aGTupQ1XRC
QSHOvcXvGpPnnKhjBJqfbnrAr8MUa3rECKzPR+AQ/YzLRGy2WkoNRcITVP/4EsTCmMjh+BUDzMlA
6H+kxGSo309sQbLkVSrqIXav1PQIpSpuU1/MJaA3NPVBSLeSBujxm1JWBtb7XQpuztZEV4QKU8jJ
mStlvEM76qjgDM08YUeEgo6bfBMAWfnpAstL6ifwmeX3voFELlW2nMjgiOyBYTw1m9aFEldNoRhE
yKkdQ38IQfF2Msn0oW8VKDqEL5TDLJXVCVyJnyWSrhPaXgo1T/o4eBphN1EVKxDiC3dcRNLxY0aS
lutPTWMR9z2l3dvlguW/LBv1ugcshkXmKxyQGXb3lsLQKv60h6R4d8wLbBbKI39Tt3Td7OSyX0mc
nL5I+Z+74cvUCNuBK9jheSYQOh4gHO4GiGDun0YNJVl8j8GJS7RmyimXhZDiyU2pD5etNaBvRXBV
gcmm/oolBOdwTKy+R2jg3xFwZm81IG6BVsgHLlx/ny9vOI+eGrFrTMeF0n7a9S1u0VmYaFYwkl1F
jQqjrPURFbWK/eSdiWezfAJrmq/PN3K97SSTvkJSSiI5Z9p8mFtu53Vyjx/huV6dKTKJA4bdE1FY
zaLZ05aZV08rbO9EbCBBVo1XfCaU6T4zQCsw/aD3iNVX7//0zVX1eneVlamYYKXQru68nFMNaNrl
3gNotCmyjVSSqy0B3U9qI9MdcHkzBVEvXdhpH6pdn6q7iimEcX0HSupkK6D42eFC3o3/UxS6kyjk
HTgdDTZRTlBwf300DPyMbIoVuvfP1Nw3sMFOtuXT/GTBlotpblsrNxvNYwF+CDYq3V0SZ+q/RdyH
Nw9CFBXJXg4geYiodkQ4aIxrMmwpKzMDjs5ayJPhqT9vxg3Dm9orwgQfPEkDNeAqlU9j8JIE/3CL
H55gIRNgSp8d1OAD3azZoauobGpYQqjZerrQ2AOyPBLTgtwVW+MKmNvvoYM+Rx0u7vHkveZ/J38L
IH90B2BpUI+Jm3I5EScoBlB97JO5cHzCDWVaN8ukZQlE3uqVQR/9t0mMI4YIQMD4ZmZ82/Kl1Vo/
EIY6O+OZdZ3Yc4Z7JN3cspTo+XUKlRj7P/Oru5R2oXSHeatoGm6NRIec12u3Gb0KlR/UulytjP28
r+qTZua5ZID+fQ3GYL0I/E/zXyt2YzLnCQ/qYWuqUd0hhYWmrAiXSneSW4lsQK/gCNMmPDSfaOrp
3u6pbQ5LGvFa+WoHPbuxDV2D0ScPD6bupKBbwxjq2oqlvCkGDSQRh2cKOzQp7GevzVO5/yWCK7Mu
/Q3jH5qI0wNiO+HpJAeyHTcrjQtPi6F0ed3j9Qk8XNhDRIbbYLqE8UD4gG8l3ag80B2SRIkYwVyY
hMLuZIW2ZZLO+LvyTLSSmFsa8UVModhZHshx4+3+vC7PFZVygN8eupnFUGToPSbq3i2jvNYjQimG
mbQhnyKqIB+2kuY+8sLclLg0rajybhm1IHuyVR91A5AQQMmxvbMmcfKuLjjlTvvucdWC5VFMDYny
K5sf9LCz4YhS1jpOZsMV33k356SA6+zz9z/UR6QgfUOwMOFLMGV2eNmBpsXReNrG3r9wXdOPEbXM
19g6KCW4Clxp3w2PtnpHJwXG56Tm49jttydZ+Fi4mU1qKMUKzG7o0EyAchYAjq5G2ALjxonp1hua
djpht8ZBwPeSVSLg88Nd0HH3P6DpkNLznpY5SGvmyjNk9eXrUlRKEtm5nVTkfzKySmcwrRiZcXzr
32Nkj4nBlPHj6y5QJ4KFb+68kXtT8XWtOQLnSKGCnef/mM/xQzZwEOKxI/GEC8y/zlgmUy9N13T0
PwM59jWpqe2+QO8ZY8gGjThptfRkj+Yb+JYt4a/JPBNRt7T9yGpLaVYqSQ/c9sGYcmyrT+Dq/7uF
vvYA4uFevxbdJTWZbFtZpuV4XHTzvpCpPeloUDk2sYNzdTbAjJYYAeCHydsZCeGLvS85v0ADo2qW
Z4kYd0lR5goQY01FZ6GAe2GZAAe+IRzrR25cJQC6vzDpN1gkL1J9FdECAwHfY8DpVet9Lc78r4hO
aoDr4NXbdcJrVYaQwhmz2c8wITVvsbqXR/TgtorTOmVGPi45zzm0IXrDn+FBVEns+PkKhVPxTS5G
JiMm8O4XhX2odgfpG4jBe7S9Spa6aKwnjDgfcE8mJ71yVHimlUalS5ekIJ46Djt9fyPmI0IYOIlK
/FwcMoVwW6L8+lbMuSuPaRHQelD8soBREFA+K6msJDGnI58Y+X9SnAoMA5o+UpSOrXUnRICdJaZT
La6rOG0OfxjdT8A99dzc37HVpRQSEwEYxPpLEcbeGzcopJdZSEgcEautsgL/m6smWpV12yHLn7r5
ByMm5gnMBEv/Q8OQSzixm+FEYoz/c7533nIfgtFVFR4JNMmG34ppcmEGAteZ1wvtkFGyKby57Z89
2ZuibuInQmYHbuHIIqQnTKWCDL+slpmqb+1PcGC1qFXCb0c8rRGFqqQAUBXcOeBmvEjMD+oFBhBP
213NTBIwajLOcZIA3R7VaPXUKjOk5HtiIB39zYE4ZymevlBniKg8ncQQJRp7NwlTnOi5hBJbV15y
OVSBZ6owMvc9KaJIWsqHXuD2KU7TpOVuuDCs/1Y5c+mtgT73VaC84BfuUDTf04a/U7wmOX/ZWrwM
aRPENQ5N0eztHucmU2xfUwmjbLAoO53M660pZNpKqzEsVXN0CaFtG54NoeZf8kBIBs6mkIMq/03l
QLPQeFyJzCTPnrI+d68pGaXSOlXOaLu+owF5ILlMqOgdAzdv4X1swursqstP5GSjOOO9ET7opEeT
SaLKW95LAJX5YPkmUSSa+J3mPyMS/YJbPHFe1Dy4TbOikDmdMN1TCCqpLhLQo8khL5TsulFP3NBW
fPqQO2EHmx63QS1tx0KSHT3Xk6tkn7jhoibKLF16iMX4qWDnLEdHF+pBGIr7AabLY5oBDiGmpKuN
F/Obr2H83ckykjK+rgKexFHPRLA0TkmJqiS9mgKQ4tREp40229aFDzypGiIxy1OIg2RBQ/uyVDTy
Dt+gHx0zzUoWG3zLkkJU0LvoUa/Pg3fU5VCKbXWTq7Pubhx0n9+4UXkJd9GdUVlvOq1MpZpTOqeM
iTNo2reA4Uc12AzzdxB4bbAWfN1Nw+QQQDciv6zxeeY0vneImaVTENjtBUItwSsfVDzIsxqU/Kmz
xz95erOBfBEULMFXpSwakKvoTaJxV1QAAxWgqZD1wGVHgiGZ+qtERIsQGY/x2C8iDspqYu/thxUk
lsCF3cjDuuhVRjYSUF5ZBGGxzo2CZv5dYnYjcuvBxMS0wDGMaLpJ+teMYXC+V7ifhMFR5b9RRT0+
S3+kqVhxgx8HCgT+GAsC9kjlEiblaq0OVBSr9GiofdsuFqRO4GgP08/Eo2G00RDxlpQCKJLpqHD3
LE3BWNJufz3NW99BO066tMu+9qdkU2psqPTEB/j5c67ufrVni/hOkomVOsqdfbmKZa6IOzrlCrQK
R1uQdHozLzMaqSSoU64ypdHXJomst8ZmUAb3c1W7jikpEkSCcRPMR3hwcxYuGLghnu5Cj6tW4K4J
LIL2SFuq4YAM6F/EukuztwiTfP5kz+LX10GqsNFbuyENdlOAw5EIH1H3yihw9HHpFC81qptaS6HM
OEBh8v98o0F/dtFZOHZcfacSz6rkztcNwFun8z2MUpQU/QjVaVTg4jUqWCPQqiUVjiBzyBCNGoCS
uAX+0oG6BoC1PKuGVaJTPvKWgY3pXuFFZwCT3LkFu+X4ARzJQNAwNpnfEhSFYLO1QIgM4aWFJio7
FCDcKSAtVcyld0dcraBQL1cc8hlZV6wSsEwrLSeIbbjUWdd5Wm/F57YUvLZptDXireb/CFB1LenZ
sio1IWguLOm/Yq5ovoWlxDGSwPU8bM1fRDdOpuxFDGrLw8NvfrfmyWJpkVEtCAcwMDmMkHudQPwh
1e//QmpdTBS1xXyFg8QAwqU9G5dt1BXcy3QcaCVMuF6R7nezlF/6sNJ0s2JYfBnCrbl3rm/+5KpX
WVdrffCgTuB7UlOXa8kRZlY+ShGJSYHPTU8dmvINGJ43NoK2xu3HJtDQ55F56ZUkFyFWef+KMd/V
gGfni0BlsIajIUOx1MvHJ/BXfppqHO7rkvUSJYmacPKsG9tFgjJluI7oiNtTeSqtnQdrimuX4327
71leVGb7vYOoDzglHXZdjgXKHluJoGz0NFJEck7veRVz3FldaiBtdll7nNe6SfdoKJV76/s/Kvw/
B38DMtG41/PelC5JGwVe7YK8F1oKnOVJKIdGhAqpjtL8/ZdEwEQIrwiaraCEmZxIZxT2Xeq0vV7X
fjeYYXWNQ74QrU9CbIRBq9UHsUaxsodJyFA3pWB5/f+7IeOgxI+8Npgp1Xfl3OJtqAxBpPXQJP1z
up0NmlWCZ1LjnaeXqX1lowHYLoAAeBr9qtCnhb1f2Cpe8Pd8mSHe4MrsZE3fMq0uwY+4Yy7c52iy
aGO9+97ZCVBV0HCQGjdECuvpu0/pmRPZNpvliHzt4WTc2rL9thn9ZiQ5Z51yoy3jIhzrngcxouAH
lIjbWYjqer2dk5JA0ENCxPAPzAK+Nx+WtGuhX3RIFCoGP8QNM57SfUzJNRYr0QRMqL/tdcrBkl8x
lhCSx0wa7peS1E0fOZSOJkMpMykMJKsYLYKp1/xJDWTKHP/roH6PE2lKWkHUxigGuql+tUoUZtdS
fEuVkI1hCwbE38s9Gue2VcINJmyhP6gTYOjkvWzXoXeBg14okWbm0cydeRLcka4jJxgfNnuLPWnl
WOa+LijGd+0k1tbtoUaZNLWi0TtR4+qVAiYwf9jxShQpmLJQCk8rjT7GrjfYY89blIRTIT1tPcwc
F67Mfc2ZKMPgqmqpxjsKrlZxhnvkBJ1Djoau/9tbfhqsKkhnw4Zl4ZmdQnvVQalbrttsRxAnr6Ht
ELgzXOeVyNuqYNj2VgdSyCm8S7q4tgDoqD+fK4PX4JNXht7QKwFzxgRCWQ74W3xmK28dftMo5yS3
e7MJtsFgHcmKSi1CwZaYAbicE/WnBqAYDuvXE55E/iNQxc/sqhhenBYgSqGEVdbjv6M8kfhewBDY
btR/Bveuouy9mlmoliCzBqvQEJ+BTnC4cqq4X8vvxAnaOBSsTIsV5Mj8LGYOsu3xTzXY5LrIUNlp
0mV9FhbCoGIm/SsUx+ghVhKYlk25Wd8GgSMz16z5pH5+v0z8lEfLFrV9nVKuimvQBCRN1M/D8VAE
4eQNTcZf3eRTdCBmcDy/fj4HzpVGBOjl4lZuFLSSvduLnGkmqfPSAAnJgomEztOvUzvRlDses0a1
MghAW8git2ffeAw+L3F6I9TtJJb4sqCoxZczlNKItrt95whihTMucs7Xf30Mvyyb8QTMZIM5F3d8
fq9sgotei9/2izvtR/OE9+Mp31x+rtgiYoEMnNS7wYqyz7MfWa3dFYjae/QHJNX5DCJFruQIvfxW
0FYtpWGIlubfomna0m+7M8sbOG7xRjR2y8mOBkTmCsFq/DGIpEvIxm/ZVKPsu2quaKyUNS08wwZ8
Uzwq/vGkyvibHotSwrOYxgV7CSWLOxYJLFcUrYf/Ob0obRtpznqvR9WMEfL4Em/6GtAkn/md/NyG
9723DHtl76ygRTJghWUaq5zfGV7DhV58gsQoHbG8S1AAg2irlTKSFg5sdhIItLCcTjRjN9Or4VMN
c7EPsMIw5yd7cK6YE1EHhuqt9XbDW+XuRaTZQGlCbEIfutGGUGXCiaiIUDkslRLWDLxuYy7hzycc
H24t0FnbSODvNiOuEx178eo/NHfWbywr3HPNFILuRHvj+JNuhhly/RwhS9hO3/or9ZLa3be6rL1s
QyODiqOrFBXC4SKUZlCanFg0RVb+hcWK5sLhVEYRjr+hhls76+EONkVlQ8YQe3vGyL6ZO2mjHNt8
a91FjcamGGSH8ysWkLwVCTX7HnRklTQH+Sn5poyP7d2cKFwlbidBBTM0HYdM9UoTjpZVJF3u43hW
G3233VMg1qZ8+DxpxQnKMf9Tc05waAoYRZ2/W0G7xEU+no4yBMayns0nIe/s35reJ8PSUKSabcpY
9j9EKVqd4BdU/SW6Qr7s1ND2qeCgPKUGgwXC2wkLahGUZ/rxait3q958Fd1bF9DbmrX59V9DPt3F
1tBVyYPmbd41KOdH8sc6rxAe5QhQvcMbJrHmDxYTmF7GOgSbtf8iaXmBLXJwSxa8DVmBNFgQwMcM
jJSYb6essiisp++ZlUO0cksc0YJPxCgFMV8JyK+lSQCbxFRfd0djYszPuKiaHvXIlbv3AsvldTcI
taQ3Mw9yDOAybVu3sSFK4SiiGAOBAjVzaS/4U0is0HIsmnHFnG+cQAws5vtnTKXH4j4w8sjAkHIY
WP2yIMUUDlzTR6/TCcXiYPbRYUIpP3u7Ow58Ii1kpLIzUCfy6hhhF9tmH/aKfAKIyxUY445cdMBa
wRhfNwesQImEODFoch8jAzx9z/xM7rBGLocyDrQqdNBOoF7cUMZE7vWaHiCbUUVVm/8yJdvo8ZE6
ssLi1TmbjYe1GiXIvh0mwWUhX3zAeBAgOFGI5/qTMFUWIhk0x7RkYILWJSBy/bUZCQZ7Dd3F2vIA
CKdpMX6Hyjuep17WKlldmL72rmhmgw56HB3Oq8hcz4m9HZ/4YLnjP+nCRtPmnNQBW+LxbQRdQD83
5Uxn42MsHYV0LF3kVY+hX2h47M/UaqN1lVLFDCJAuDGBppyhNyQ7W1qspCZmnIJLTJlFSVINc3Mg
HGO4JqH6ifD/8D0JiZW9ASRJt2yv7hG0qsBYe8PabUktnCBCV7CRoV/lUoIeiYZXuKIvvjlrwUjE
2G+SKTglae8tZob4OEamcZE9vYOMhtJu7NL0J3C1cHO5AM+7128z+LMuElyKrxUCjVcYp2YtRBKz
WEjAjRe44+d1GV2h1Fi6JObPAcw0h3Dww729ZlVjmNzhlSaFzVPx+8TsK7YfALfVg1Er1UHrkaeU
szodPv5CBW7JR8TA4x3X2iPQZ0Pcd+X/TURwPG2t7JSQVpUFqmkFYtyPhxzvMhhrjqjEOrkWUP50
Sg40FyCCAoY+nu01GdwKeSWao2ACfYS7oXGFFlE+qeAl17XFl0LjaFMhPURYlFQOfWMAQruPFe9Y
TuHXq3fas0cI67fl9mR1OFV3+Bc7zLjLSwS9CDJh2VDq4G/7RIEWhV+I66/AikVf9q3TOQNqZq1u
8Gc5wKi3cC23UsnBaw2Pyfn3w6TzGmSA1dX+8U9G5OLKOrtdUsLZYqLhWYQJJR6JBbFFYLlPSFH/
CRxyrL0eR7AeLULQnyWmNTPpXQme/QKhA++deDts+/NZX7Ymeepx/syVzYwltmLpdgzI6Fpa7LUv
xDwikz16fh0MA4XlClPePGlAAf7pZXiCpWkJBX/dmStrfMs8BhvMCHEDOnGbQ9HiazD35ym3L5hh
NAfMOfFX66rmCKjpIo14hIOuzMeVep2MY/taPk23bXkqdsyJeGOXPoORyCSNy2SqlHcWEI78Tvkj
RlOhvIllK+CaYCDusw6WiSOuLNllW1WBKfKYq9PfIg1hieNOoCJHR8xIwpVvtnBAPWIabIdogOEv
T6jmztUpPRtV+AfvGK2hazQbeLsPgvDUAbEj2thGqEAmguj8tcYnf9BSvS5qTGPX9Na99RvM67/D
H/dID/bM467LZvPhL9zT48Almo/J82iF/2u/foJySQSpQ4hdq6AFl3tR/dhxsWxsvm56Tnf8PgmO
Cy+mQqO69fJHP/tsZoHN5Cpt4ii6zjlIj2xhDUAHeG2g4Kl7rB0qb4QpwyL2Wl3TFVewLIWgPSpU
G7cHE9Tv85sXAUdc7ziqrsRcS6FJ+wszcK0UjVr0j2GmeSH+lD0xrCQnJF3IIm177NWklQUGxfPi
6uoCZCdEjdhP8c1ZMboJMkIFB3TDnOyrlyY1Fz1C+leZGv4YPzamLs2yHttiz5EOU2dl24WVrF/c
g56bTjOJzLIaPYfrI7ONz0BkHq5VX22Nw5tf6LGF+v2ZTAFBrtZLQOUwRvWfHwy+oLuXfDYyblHb
DyMyXYTs0aua+rFEtr3wi6wW0OFD1DLqE50iOeMTk+bWNSjD87OyMGzBixTcgFYgjvYs1EphEkqC
RYaPY7kQZI+hDmaGgYx4MqQaCwYgoM3p1luDWxmOnqJH9R0qWSfHgaTW98SgPR1c5NujTXhWXnNn
dBtrDbQbU1FP5kvN3lt7kUex2TMHx4N/9e2aAi/LGoqh5gD/UBKkS0OaGsJbkOPWhHXLC1xEkP1q
Yc6WGQ26Skz/AGhoNWfBdacU8SPu+R4ugsrXp9abvgwLbKNSArnKujkEEk5hTJlW8suEHWYfT+m1
uPoqf6+X9yV+xetnS6EzemYJJ91YseIC78RADM5wDj6Y4ZGwbANPM7GgY0xMo8nEq9hWhzlrvW/J
xFwhakGyh4Ng6TmQjoP+2MNZ6xtUBXoV/8XCCMJM5RyqE5/KV4EHPhnzPFxJPxmLQ/fN0DgGK+Oo
v60WBH5sEwBPkn5wxe3Sga+bhhPK17Sfd5BFCPnJNu7O+00BppRJ6xcDyVuWDa3tQuq6bUbBhNrW
44psgvgdAfoT0mvN+1Qs47Z1BeL4A6+c1SaAoAbWRLQ/aaBenWWqxQE8HAfmQXJIaSIM1Heb6wxK
WraxkFS+p26qUnHTpzfztrCjR7vqJ4SQt6256hVfbLVYuGFjKHUTtXPgGUazFvm9Ozn250DQLJi8
3y/sHTT52Mnq0FUnqkNLn31RjSAJOnd1MPeILfjr1a8euH6PsThtLh2JqlpJdkH1oKK91+FKM8Nk
QnhsAl4X8D/i0m2brJfJG6ORkV+AQwtz2fwVmVDmE3o7CdXfscIJ8pqf+XI9yeATvAi97wVQglrg
3rggG5Ol/3PoL0nP/gIK/nuHzJsfoYwBzm8bwRUc7kIgrVz+JktW0DLRUeMTaY8T1+jHVmnRQMb+
PHUCzDUZ5rxmDXCgpPXOPPwvd3KFu4dKw2pORCktFuUTGMbHhOwm0OxYXT0gelYgE0wxAv5EFgrj
ZJg0ZGUbsGgwkUjKAmwK6mRSJzSmdgeQyJabETvcjBjN5E4+TkOHP8Vzn77ieHdlDPamRxRyLBwJ
0V7kZu5/mZOfODg0zY6MvdTEv2I2kKni6QvWDrZa0aioWyAgDnTzR40UdKNJ6RT9exDwdowNH86Y
nRFwq6/fKWkqKymrE+TQ/2deYwINzXOyTdcCJznBfpClejmuvuIpEAZ6pIxTlH+klFYVL1YI+nDr
SHQtG3o2wH7utGVtKWp87xUwo6vDvYJR+x9g7/Ecgc4HP/9lzw7XghhbigAlsKHTOtzjQmXspyll
xcTnEXWHWYs7T42NmQUMASA+YSFHd2Lay/yAmA0OzL/p9FBazjedde5umkintUd4wlFCZIQ/hOkM
haGa3i3pYUeD7f8u69pWvDnZySEar57t6/hlsiE/7K8EsVpFuCra4pA78Dr1x1yjyhtFYzlxqheQ
JowCqFHV6DopDMfqnOY/lR0EAqvc09iNeYiC46+u4lQCkd4PO69sUdbEo+VGF/6q9g8ZMVscKKLY
2fq71ym6C/u5mGdUgdFftSYGQpBaYqh4pnEVBbcaVlzV/wlAa8yXOJ8+hzsUMd9I7ls7ndJqVdtw
ImItp+NpJ4FMSYDjNe0TDJXsq5NUg2rtDg24rCkerAonhX23L18V26LlV2lYvhgWOWNPeoYBcRHf
T9QO7ZhTH6Mn2d9bNnQM0z2AqUyewwmRGZUtUNQcIMQ2Z2yKkqA2vhZv+crAFECh9pYt5+XC3rzk
0fC5Ci0ON540b6jyUtIxy72qeSZpbX0rmOAP6CeT3Y72CwGp+dVqHZB16+aPVULvyvPjF42xDmJw
WSZfCFCrCxAjLl8u7jt4Z5SP7XCHIM8tO95v8n6jWPTAoAUKQReoyv3+NtmbRoS6mGn+zbO4SssJ
0g0kj3KsOfwHal3Njh3M6fVH7ay3jae5jweoqryMv1AuVR5ij0Gnys9esw7+sb/JNeBAcUtanRZp
WtwMi9SDXqpazuoRVGpx5SJvA7850e76N3n6mTKO0vD1fOygRtAN2Zcb5vkjeda64I2Luvrx+mUP
EkfmaFu3Ggjs3UnK4lVoBKXJRc/6J+Mu4ubomvvm7AFG9hV8qd9gAKD95kmZ7GyMNmNe7A7bJ1yS
lIB+pRfdRg90DV1QAPR751y4/ywGV+qNensfB4JCmpwSVzUxGFbQm+1ErYBx3iCidGaCTsFWezXq
ifKjSCw6zAG5dGWZrRj8pRpOs7TG0zSPqgZxhCWLNm2SoiWEuPcyREcqBkwk2Cy3oz681AeqFoo2
ThWoEkgbp/xDwvubqzxt5eqTqKo3EKZnnov4RDAujGt/VM5z/Cs0tWrtRIEE8xjDftdBSPJ5kXdm
YkDV0kHi+xgBWwjmGbeITok9u215nXAtSFm7to3jIkL3YIDYYvFTnKz0oBFSy7hyzdp1Nz0rWhC4
5kNmGFQ7cUyLfXm5HobSDnj15m5urfqBth4yiwKPpB5txgWyNQRd+1tAfq+pWMGignz9DgnP0KFg
24eclyjFYnp01skwOZFw+BVXiFpqlFvQ5cHwSwC+Dehd/NpQVw6/R8zN0pJYSztzzY1V0XuHulI6
bcNbXP18p6n2wxm+iu4xxrpVXgspCliukhmAVPGgNXERTG9l10+3AJNsp+V08Tk4jNdZ6NBAi2z2
wmeGuMJyrkxr8MpXt2rBDvAsDGLXHiWp5ASuibqw1hgDOlNnQl8a/8+Nq4f1NdwrHlDMoTzLSK6S
eEaxthUKub7yusslAoMQhPYIzQxLymTZftsTvyI0zu7TkqJYcwwIBuZEwg22NKcHa37JFsE1jc+y
bPIBFBpGPXe1L2lj9zxCOsr3wPh+o4QSc3A2Y3jEGB9a4Tmbbx4UTrZnFvfPtl6K38N43gThJc86
XMguR/0YgX5Q5DOKRQFTaHZQY+PZrgD9FXwQTUF5E/aXqu5zWj8OCTcOQGpKS4jxKeVz5jRfdxZD
xIk5qWZj3Lw9R1s9YXB67JFn49QOfuZND4uASQs1S7ScjUe+dzYnSXvKJuqssXI+0JQc/AS+ND7F
B+uxPLPEYgoebDL6xDM2WgE5eq6t2bg0Cy4K+4dqkvxmziRI2rYgRb1xAxNX246RX5fHdVJeDQbx
cmVzkMFXSFBLnTQse6D4f6bwPAqvla2HcE+xfsVRLedvW83hQZUOJp3znztvZgWSgwbO2Ccq8EuR
9gYWfTrGtlKGRQwEYCG3jqvAn8m1SUFcHxE8T+dwOk9SEAqFdHYkuy7ULtX+g4JAnfKMuq11Ucp1
0AMN9XsuyYN/xKOaP9Is08gMg71Mt+NzH282wtkl/uKQs3urNeNc7egSiXC9c0sOhq5eElbg3Tb+
0sdstYi6fCkP4mF+X//w/jGxAy5cDde9q63e4LAuFyy8OgWy4xFbjldismkKO7XY11qH8D4lz/Se
dD3MZOoJP1DANCmcFasCWpxgMUAUsBHg2YR5JZtH69zHYoIfsz1pdaaAuK5agh1LTqb5+x69GQ9m
4lbxcD0+GLakJUZxA56NIOml/+wdY5FLU7LjFU7UdVvDEsen4jaboulZOP/slQasESaCBfm5tipJ
JGNmVoXxqmbmGWfv1oq23eIAkyeB4tkuZWOg9+Sfk8ZfjJ4/CJflCjyCbXtEWVaICiwq1NfOKrFr
JCvqtn/laFMfEbxEV76SBMJC9k1s89nqurzi4IAfGwV7clKoLds1sgzVX2VSTT5+427Iw/aHBhJs
DUL1hQIvXsbykNnLHxrQFGgJu/kedgQI8kHIqJczNPS2PFIWMRDJsj3twxN4g4QCe4ByRvL2XwIp
z3A2RpLR9dsbl2pN4k2uYjdaadGk2ClD8zT+LP8zprtwT3pXimoZVMH2XJNoIZcgBxT0vVFhUsfC
GOCAylTX/rc8p4Rh6u0xY0XqwHEGrn8iS6rm2+H2fQXo7mRogby9Xy7/Y7sHHPqvo5PSyQ+Uo8vr
SuyfCMUIWK/SezA/4721NIif/0gX7kX8jk11bm0h1hFth7HQqjjYtlAI4D/dcUEPHiJaf/9vjUv4
kUsxvwyxaaYcC9ljd5h+26hOsoAKwsji93PbvcqTka14xSjlzNwAiTbP1zgiiOMesFmQ7nXIeEoh
AZxW1SSCYWyNg1taWYh0FNfU9YCGMRdLq/uwPX3Qm3yU/P8f/BZ2OSWplvjRxWXjGg40sa0qSnBC
APQKOEYAsfURLJ17clbk+9EsRQayDubmZA4T8xcSVeTOHUP9oxE3KoKr2vaTkG07ihmAlFOrPZ/J
O+Mowv3KcEUfhpnqnc82L2/USz2G6TPQx55lB/xCXYJjvUYZs1XSjDhGqaYGvOV8QkBH2LMgp2+X
+l5Y8kjPYTWf0HCQZ/ne+te69bt+YeoLawCj6SxFhiEhQ9C0RmFG/SzPQ1sUpCGe59gyrWAzmWkg
ADmMXa8HyGoPdGSZtVCUibMjsJlQe3nvbgkkQkRw9S3hZq1t5aRjGykJ2zKBGDr46tfVOEX6gmek
3aLHRyfH+iPM+c4gPiBxfIQNrJM6PKuR6fRIPywseiqRgs7jJDWhPWEQbIJAiAlIh+/qaiK0IFzC
IEuILai+BK5b9N3L1jm9o/vA9pnGiIOTIwJPYxS07GGXHZggrI56O0BMY54+zOL7bfH8dMgXyyD4
xy3J1wsHA4FmwH5GzksWzsDkkBLaUWsuifIeDbiF70UQvsZndxcg3M6/tNkGVJ8tAjnkbnSip0tp
YBNPVV4Io5m75if0JBiKFYFQFVn+H435iAYXQoHyXWMmpgQ4RqoOttmjOXaNxox7CZAVrTFptTj0
a1x5MadDIrDSA1dryje1OPN5GpTLu/ZAdWd29DuhS0H/ofR5C3eiEAdQl148DUcQQ5NyqVqbZ4i4
XazryVEKbTUX3BQgxtDEtfN/2sKCkRGdEBK8gJa2LF1m4M8Fhv096RL/qzvsGwYxTg7BVz8Ij0/p
r7SdOtEZ8WBuQKCpuYX3ePG1i0D41xFRGjmfQl19/vwKOsX6x19ddrs718rXn5uAfdepVupfU66B
ON9pp/sNbgEzBtNorQZ9jnLrPkFsi1L+ZQgVZczkwHRlacXlxPfxKwXsGIufdCV7kYLFAFjJWiV5
ZVagInfN4aW7GF2mtzNWCl5gBw8yxf3eckZrPKeim73VAE2IDBRjnaVeAFiPZi24FVShpPMJfwY9
JWORbtzcW1MYMfHDVSSw0/EjpmTynZJJyPTyW7N9x3O9mP35Kix6XI+yNtY+kdLqSdIfFRTZHfuT
uHM3vJXbhKYYheU+f0km2YbCmKEhSYZgXurxRRjVVGal6yeajPTFLE8VsEEJXaBOkjzsWo1s5MVS
hVhwbS9FFV1cyuD1cZUpjHudnMhh16ITFAJh7//kMCTvdb2LCjKz9q+wE2njSxkX/ZYLClBjWdr3
Lv+IJOlO1FIhXqcKmX779gJH88bHUTkS2kv6nmCiQ3stcqYzHvqdW2sTO6IH1ebM72ql1HYPQgfE
1YpoY0B3u6OGKkBX2Lc0KIH58nET/V7VNxfOQe8tRDS3jxf8IdI+yIUuBEgMdZgjk/BHZtxAK0+E
D+JKOMTvzL82h4+2/cOJP8my8kFdwjz9p33oR3g/H4q/6bkc8E/VWrLnuCX4Ju67Iu4I06DB6H+/
O6yEtmViSGTfUyf8AG+cOgxpZ4M9sTVlEsg4RN39XtRoVRRLH6ldmVwJfNexvsKnduH+AWUO2nII
+2BwIl0Cwu3N3EXFZcbypCdHoGeZoVux6YlmkwkW+waRioDSdMpJGx5UN+CPsI/TuewL5ti5BNkR
2gq7RdRTBX7AerOlvtceERDczmZnqJ1Q52YMg28ZgjTQIMTMnSjRdjh5FUHUtKlRybO3jGsk70rW
3mZtVrVmOw9bFYF5pyFdVlKvlfizzq6DIvrVkygDgJqgZAS6uJRonqY5kL1JpAp/QdOc28W0Ue24
icq+3Fij4qok1iszGb91N2iS1lzw6K9qdr2Wq7MstWmNW8/7Lrxg7HQ2hpuwlGmnc5flfnZlGOhz
CwP/DwjRjvt/bgOlLPt9lEjgUvAoHNZ3JpSqOqcG3zjzY2cqJJwCtGmXePnNl3qhmPO8nAD/NzN0
fVCF3odXEKvcvlTiIUSF+YwvBXMCbEjHQPV/DU6OwErw8GRqFSJVpjv81GL0hapLeYXF/JkSmcbn
uv/PVVvbk4d7sFyrOoB76NBEsY+6aA/D+MspNWZif+6DMk6fKt7kpoP6l2MtFKCVAuEZVmXZ2i6e
CtzUTi4z6fiRx8kPnVEgybgNo8XHs5fvrlvkiFd8ySPbp4Hxm6pDVETSDVzXeub3LBBwTbzZwLI/
1ZLhuF1PMc6qiAaU2DYeqpSoNUNLTITrVRNdIIxlyEAbwlmgAYjgTYABf3MCQF9K11b9XOZgJMGK
GvME8ZdEjVSPES735Tm+nELSWIAIikVv/wzEmX+DvxiaOzfa5Abl+xt2ybYci52tdZeDRwj6QpZL
ELy4h6i3Xfh2aiD4tWlS0otmmutGZOWWtoxtx9abQBdh/WofcxPocTjxldrUD4BbQbO/xpH0M7va
TpXGkgvwPFno37Z0OWXuD8it1szKmKn8mz6M7vXlssLwyRjGj8Dprt32kYgxYVWxS/T3GF4XVKj0
89G03xyz7Iw9kk8hhFUe0XQYV+rt10iBRNJtDDu0+M0CCYDXlm4FX9FUiRb+Vk1u2iHPuRzUdvfq
evX820QMtdjo3XGPLS+y0+EV9GkOqiTqcnqyO9ysfkMxVhbgp4Iyc0JlQKx7E13CpD8bUGZVlU3N
9+cyo7F+nj/f7zK9ioKb21ZGY/EkFXg9DpinTBDNy2S/Tfi/QNWxtz362o6uLapkMO6/bNWoi8Q+
3IYsYvkBepi21efCTmzcbb5iylDKZm06sW1afesPhEAEhWaxZpomKVjh1JES/PgHX/HG8aPnPAPB
bA/gSUk3YA6zIywDgX/A+CWAT2VXsS23wWLiHO0i8uNVwnNc4EWCc8H1nKN52LyUeu0agO7QVueO
R1j+XQNOrXbxr994XuIgoz3fGhtlwSFdAbLlpQgsAki5zH4c5TLt0IDUvmr0gnoxX0ppJ7NPJjbP
4gZ5rwzdeIKLXbS6JUdTUyaAh90PfxMniPSh2fIxWTsQTfPQyD15OeRB3wShv0aBWNtusZgQexG2
BrHBVVImqhSkSNsl6hfN3BTyPui/8D1t3I8hvRo/p8UDDwoTr93HVfEPLOGG7AuGb2RJtVCOv1u3
h16+XoJ5N8IPcykytawUdAFN83CV5O7paAWODzyd+vKrwSVecN0hfYge0e7ailbQPjQJX+f8YY00
NKA45N81QesFviB6j7hSE9BaF2u3FAHks276Rai/rAqrcwGQRUsUFna+C5ra3NHekJGRQs1PY4TR
D3gOkdX/f/Norj5mu5bHZZ7uO86dgI5BLZjl16DA2Hp3mLCkJtmkc9AmzMFpyXBxJBBOsA2mlDW8
Fzp308Axf4i+pG7MP/YZc72lE/0hUPI6bRw+8q9nqZlptZ0O4gPey29Aquva3PvQ+DPggsilqW2h
4ZMIlK9HTyYaRRBw5tuTUV9iwqHdxqbsmxwIi3R9RorGTkUctBiFBu7Ugwb6Gs8K/YmpKh6ISiJa
6igc0iQcrHg20Rs3mXNCH/4/YU9cmCwLmkg3C48+vkHiahn5aE/1AL89+el2T57XWDEPOT7hDzz4
pU06HxJEcwmLpZrNocInOLsRrQp+No64cCk6qwfA913ngGbcst+qaxoVGlTj+ohYof6jrztUWZy2
BJB7fsYhmrdhILQtzQyeDUBBxSdq/eK3mgQLumWkTukbilELSY7e77Di31xo6e2LNurqKnDOhOCn
r7E1Zdb1b4IRQu7icjmPUJifaWNNk1v7WSuz6QT06BF5rdAe4WfuBUWBPJXYEE361DhrElL/+op9
WLWpea/VdCOh+fu73m112s0eulyWcHobs4wByl4mmSWfIWum8raIvuLbFc/A1/tPgzevHMei3Yxm
6mgMkINF9TREyGLkRmgTUqMuGxBIAjlojj4+o9a/7O8oAsVMKZmwftGWRdiscMPoPS4vPWGrjsid
UXaOmogK8t0Gg0D0Pu1N20vS1TftRiGteeXa93eYiXt1PLEZv5ERQZzdSFy4hu07qSCmuHjtDXwi
jKoTaBNixCH/l1H4lPpDAitW2iCclbRegYZv1zv6oq+9imEXo1NXXzYCdMuVKlQ4Yi8hdKIkKUiW
ipIVu62THmnfXVhspNHqRAYPKmkc5sv1t+5yrc7gZEPsQewRK5ggMxfZD2jwp4H5gCWZCwkv6/2F
X4KK4uTvzEKZPUMiVmz/mK2h3leNqKh4e3dHmzJHB2JukHnbYq2v9mQEWhAgNAN9tjDlMyceiiHr
B2ohZiPo1eNPYRLv8F4ejvelIHh8ZNfT1Z7+rY0wu9RvzNZh/JspcHzRxEKI8CGMVCnkVh0YKY8Z
Hkblx7Q3O9ZgiPApboBfwlKYkLEjwNB+aO2535tsSj6B7Dc5XzUxj+MA5ATIixhpgl6cJwnfPDQ4
PyIt3zpqy94Qz1aT08Vs/s0yvtPYO8E6u+xPTyXtF6/NPg9HrBn0zsXMCu24ApgCpeGVFz8OpArO
tuSoyC/ZLfqUlETcqm4qyFHs88UfrvOnMx50E18X9fQgJd9Dm3NXqKIEXy53lCRxEXpkQ0NgRnSZ
hmA7jTelu/YtFw7OydEicHl5fB+Tj7otzruZjDwBO03NvqdklNf9ybL97+48SrWfnVAFGRTL0+jU
un6oELwYwrLd6QC6gb8NcNJPmij1Ej8dpoRuDSPoMOLYKVM5PO2vmuc6P1FwoWegHUTEFCz+DVfC
drU2hbppoKzTSZ747plHgeqkdRYffmYDQRf9hFZYtAesHDdmVeBPG/7zgVsYVMkPb1LXW3pfQDCC
0jlKJ7P2gW0o1s/yQgTR4Imzg3HSTgB5LmID/AcVvoAX0TR6mVGoJ+IGOzVtNxJnuB+d5G1t1ION
LEUQjv/1r41r3M2jAHhVBSiBWKCoRe9gs+YEA51B54nKh5o/Lc2wdPTb/L8AJzJJiye0I4/QJieo
DBcLlAd3AKWnTa2r9pOXROPRhbzCF6OrYmtd6gJYquKVIrBStPKwpvsAde7qJTnj0PwN3a+kspfq
kYmQMaJfQL5m32fI82+PaXdTVRepWFkvM370UbDs8pnhlijsFpl1LwOqZq1Il+Bpr0uRBjXRWlAn
JU1Z2r3ezoDZA8K/W6Oc3BdJTJ86MuDGDLdF7j5+aoRttqtWg81JIqyFco3SEQ3pNZg+j3ZKwwzA
gDO5UJm8uL34Rwjtw8GlNf+kAtXramVbNJZZQJd/+CC1HL6Ossu4K79ETiIg976R2K5xjikUOlpJ
Ubb1GPsRuIqfynX8RlIsv8QQs3qSzT4+kIg2J35ZTHbFBYUrvwi6GRttzVAMpQhv/htjWOEf0E5y
PorpTV1DyZuCdHa3wiQQpwJ9PBezOWCbwmR9su4xwC/sKqQXbpe2EP49PNBizZPPvRQKIjShZmTH
G4rf+inZz7BZp1/9Y6CVENRO4wt/Mrti2uYvwWozrRWqN2XZfBYwKEg7R6WiMYp2jk/dnYOhqrlz
65S56GFDsU5haTO404TaXso+3iTZBq09wxSJBUq+BEIesRNUZa72S6yKAPUkRoipAdJ0DiJENGHu
U42yJR21hPXxzj2pI9BntEXeEoP7MiCYqNW/mX/oMIZoy4m/PlZleFfJ/U15KPguv7bF9ycI5IiG
UEOusil3Yo+WpnsfoRoQrZqnvvqR5D5pJml39nft6RmPD6p27lYRDdeqztFJIqV6rLtO2vL92+Hx
wQHRd7Bw4ECO1ddeRtUWTRDM7RSChffyoG/qvRsvfg/VVIprdtDml1+GqEhLJ/GaAQTE7osRp68G
dy3MaNrejRyt0d+W54p/n0R2+q2YdDua3Q05gmkCFi/OCgvW7oGqSOS0BD7hAffcEyDPQDkkwELB
xJBSCU1b6XD3zC6LsTQg+O+WIByvxvu0V8EsEGHN5jiHGRWfYmndh1hbzfktJYQK+1pGNMFZTQPy
cDEY1PZF6eocW0LTLSxj2SacFAfk0aR4/qpQaT6sJcnHj8pMl5Clx/VtnWVNKp1gz5L23ZiaDil9
+6z1YG3fzpLBtf2JAPkpYZsZAmoWazFvYABbY4pRsl0LrkVnNQrMi/CZVmpWC5lSrQYGsrmDettC
NnY4ZwI7yEz3J/8zpij77eT5Bm5YPcBdxvTDQ9q1a2NFdZdJjw7iI0wisGT2WfsSBj7qmg3XKZtR
fEWRAFws5oxoC22trO4lz/I28Oq30zI44nI+DVSQHqcKROOclhoOyW6EbWyDsql8ifytA3CX5H+3
H2ywcOzKSRONtTwZePCBQGk7Mwa4Unsj3cyUH0HZsl/BAAMRom0BPf8nna1S1ftkCngcyuHW623G
c1gjS4qaJc0/5LcEmfPbSPibvuRwft1iP0Toal+oQ5RVJwiSJN4S4DHZF/47zCG/XpxozoK81dX6
02IMGdXDVx9DGEcTd4d8YofIet5V42D//ETgloPurDJaTvK9G7Wo3S7CX+keLGn0l02N8Ihx1npT
/OaH3BcbgmtFu0PLzF7rf+GdBVW5MEC/NRNFVrHcgsROzOvcDShYEDNbwRX7M6oFMcnjjS+3KZia
UMZXcZ5HNg4Jsue2u2gYEWeBk88fLeVVMzGzPgx+4mw0qfZEAU28YvdJ3A0vFk1dewfRCBFGq6yj
DmPgLKEcP33h98TPaz+3z7133Kk4uMVeAnfnaXn5jSxv9EJ6z9aCK4GuE8wJqr8R1uuz16CMKQ8r
azcrmeKFSUtqn3Sd6YbziRyi/dn2/1CYShc+BcEw9FtAs5PMOJUj9XP4iT5yIWMD8uw7vpz4jG4S
nuvx9S4+B0VSR8WnajZXXrOtjRDz+2qPzVk6T3qIQoeomRcYYReBxN5yOu8blfJKOrW4wfgDR1gB
nvqOSklURj7cKDSwi8txmV5a0Y2rgsSf5PCu+NdG42dC2hf2mDV3lA7rx8Xo05UtImOK9CLRlGPn
z6cSs9j9+7G+LRq5F1B8hfta5t1qKMYf4JaJLbqutinAPz60zwc4KOi23AUFRK4CgQvN3WWbQrnp
FJU83NzdOkfSnftPROiRE0JqKhBffTTB/eShRH7qQRAwWPhY+S/PN8zJKWC894BChI1KlUE+QxCX
S1kqDSi25UJrNfa7Y8q2HJYf3q+bAr0ZH0lAk6fBtISR2AShsR0occ/63F9qLaoXYzhZBEo2BrsJ
ice8aUAiC0CpPGu0HGnYzJ/iSavfWtoM1H8Ud6MBzzjrODRGA8jwAciNuAiSu4xkoeEr/vX9QJq/
7MwFXdBl/+DF9aZVI3JNqvPL+/poQPmJ6+aTEo4FZ4wTngQemw3MD+C5q7ZK7FYTtHoUiV79r6gV
jyC1Y4krXxQKJ3W6F3P0Bs5Te3YqGu1ylwWs1SB/Ddd94sjM58SJNcJGLSzdzjPpRcWfl1NRkUa2
ojMIw0NB7LUCYja2nY8FyruZM4uWf8Uhg1pKDayyUC3q/ZKAEQLQXpfi1zHm+7mCpFD7s0V5To3O
rU9kEWUpvWdU3XeoalO8cKKfLZxPgMJSZFamIh/vTZBi0S1NlkOUu0H3b+4gon59NkFqGtJ9WWuf
WAimG08z9CeFQfiY/Z5QHI1uXNJ/9eHEZekQGuOkY92jn1KBjwUkD+TTeqOADPnZyVB2QGd5IikN
z7Y1c1OMgS5cHDQocpXyuQnJ6AVKyLFXjwqOa1tlk3Szer+KKb6Y186S+VXkMkcfLVsXi/g8aXdi
B+Ao6vDUUqvidKpujyHfvMf4XZBYI0z8k68DAwICe1m2XsIMgaR05bB9vbR5AbMnJ1nzE8yV80yB
jnutmaiFnhXbTLhRu15JRiuZLbRJWNEFeIEvH+7mY2w2YwZWyqRbd4f/UiK5PcFolvI3Td3lrJ3w
w3osu6ySJaoZMO7xtP0OHC4bSupvCLoAkn2H5Qg88v06gX2Gy0P5nH93Ae/pcvAHwBf4WFsjKP29
lAt2bdTuo0b+MD2HKycAfRwkLSzxVsbt3i0WkPlfUV76ryW6x9gPcDX7lj9ZzSR+MAEKd6eI5Y5J
rudaPSp5CSWop92AZCoUyEIdBhCNJ6KTQB8T4bvUIVo/MobrVIujPRQW7n0H9Gk6S+1N7v7eTNG+
SGkJebe3el6ofNl0V/sTBd/0H1zcezlPvlqrKMeO1xsQ+Gag/bgA5/+aim1csqGoMRSfFyHxaKcD
fW2RqNH1OSih0Z8D1A310JqBXoZHcA8WqSSwwjs58t0mjkg3PDh1W7PwEELboaNlTOP40c8uUep3
3/kddW3zChwoTbFTb7XBExZUA44R8JiNiFsLt+et6jSNUIHdrAtP8xNE+9TDuVdXsSPNUtPl36gY
C3apkZEULRKSCSKd3ZPNBYJ0yYVGTSR4fWC+sOISocJzGkko0VsUjHvuTSm/HVWJWapb2vb6xme8
M1ycGYZrgHQoqvQWxeOBzM0+2ZLkUzGpL0WH73FiLLJBEUsiRGYpiJx0yUtsHCZsaYpzJ/mqUOUH
Pwyl2nLxfGUcbqaj1a/dJc9ZQsN+zww7cC0ig+ErfBpMdW+D80qcVJIoFS4ynKX1krnPcxwFui9M
6ccdg+y+nWbkynW/BjhZpC0bU4vHXDlFZQAiFIfuhqIdTj8zGlMrEDevppsqKgXufdPjfgwib07e
xlfTwhJOuPCJnR0xVQi669r4ZWVlVJNMcQgGnoswcVAVpq3RCCmg1fzKPsytWc+0EkM6Ywr7lcYp
lPLSKXDAZhnqRXSQWpYBJQrf/tM/vpT8I3olwz2mghrakTdryMclOv8bPfDQyqVycbCo+S/h/t9p
25Pf+Kueu6DsqTo6xvO9ngdAdAU+MxV/wkhgMwzSB9CC1Fuk7Yrz6TPAwSySw+JUsu/Id0bitGKx
ppFqfLkg41nRKFaml7FSgvNfujW36jcx+miZLNgSNagH/XvHkrbZf7+NYdn9hUY12Zqrs+OeBQ3/
rbxXalEjssay24WKDBIQev3NuPf5QWs2GbbEim5QnWhoK/Md1x8baqn4OJxjGpKTqJZWlg57eZyo
vF6Rg/uRwekQDhEvPz5sKU43QdHfavtIkBcUEMGLqEtiIIpd3C4EUb+ww9bNTDsqYhFE5j5qHuCd
AMLvkpOub30TusIIlTG+522Fa30xpvipPQk4/0pJAev/lBPOJgalU0e1uANrnJ9YLRA30YZJ3LRl
vRq6LM0JvBi7eKx3TbnbC2Nh6H3vGDS0eE1d9aLL63I4Qm773FvpWuIOapnrtlTDJX2L7l4jYFft
4NHezr/rM+0+XmG6PHbjtAFwWohbQ5kXBop1EAB48PPMJihJqMa/OKWBJW4xaZYn2oZZualDGzWm
XF+6SDYJgtGVSPehPyvcO/wyPmiPNY3704PNI2uGGW8pdAvg8WF99qm9QEx8vvxrpbf3DgHE71NY
jx6jwvhjJtg0etqRlrJU+1234kB5C/EbRguwctE1+SKKE36dbYGF/THNpHTQAJbXA2Hooy5g30Hh
wUim7zQTDbOIMfL2XeDX5vn5mND3RrCq8tQuMeHsJpvzq69tAMiQpCcr67Ou4zE5zzMGkmTnnmjQ
m1IuAmTwFuRtSa96Wlm+T+PWk5qwzGXQDXUJ3JdDaY5kbGGRbqNtG3mrfboYy+1Al78ZnSojJ+Qa
NCfQ9Qj4T6ztA1ZhP03xbVPnTc5jrtgWao+WhjN2v6GN8lA7DIcuR44ewBgNDNlTAyuzvxfQ5X/T
OFrWUs73vsGG6hm9qqju7WC1Dk2Nq8hhnv1g0AAsWQG5QRGzvYkwYPWL3aBMv01VofEVevDUovEU
ZdVq9Abbd0z+VNVoeg0fL07Telz/nFjZLAvQ8JOUNQzcQmetIvajDbsP9qTIIxyQadb2Cnz00cwn
IFm3y4eBGHzd1LZMvzEhhu2e18AvSZqAPCwrKhd/sLaMn/Tg5m29tcUMhOzIqIt74NHdOdH3/k2k
YsxCHQmFLW/mMEObpOdWatv6yDnczZHyxRqFRzzDHvDAuI/Sea5dsyR4iS36WeXGBA6YC8ePBBPj
bMFgbcSR/MeqJFJLXjPXgAyUdjLC/EffjHZhZiRAVhzFZH77zCQYyEmcjdw5yf9snANTZbjnvpjD
FmnXWgJE+7RoZmjH00AXgGfUwCwsGGvrz8+C/kVnasmklj36Ty4Sq26pbAcG/cdckDVBDznkY2DN
QCIpOmCFhut0209JEJOgVNaa412sUrpQ2dd1v/JvJcRYTafdpsJg9YbanEGaXvBpxfYMV0WyKfyM
bXjLJTtVZ2q+woohpSkhMoQhCEXv4RBt1YcMLb7QahCyM/CcNK36cv+Bk28TZKi6C7glr5RIHxiL
1QTKrO1bC9/2p6JduJ9OLgGY+BnqrGJ1cQ1KqFHtz692xmtUFRsDC9UYm0oAZRHVcYswORl2T93I
y/g328dZza30igLLnwH/LlI6K5cra6EvxCF4boIJCqXIEhhoFa4UzuqZnGZ0rQw2E19KscK0zgjc
vC7C3X4kYPrd+9Uj4ctJ2sX/JlzeN8H3KYaFOGgwHqtolowOpu9+Bhqj4hNRIRnXXyfoRsxzSE6m
tCZUcCwBPWkZ4FB8nwbWzWo9NoWHUC2WuTv1RSbm713c/WaTokMYdKuR+PFZ398Z0awfeaLkCuEx
NPqTSzak56fiNIvIm3ktMdHrH/Yr7AltxryTNIqt5f/AZmTbZBGj4aPWnTDJBWXItm8aIvTCG8vT
Kdy36Kh9ff4Mw5fu9fyhzagTgjuIoNNiGUpZnsy4mz101Qnz7xG2j5eQ7EnTRyQDA+FeGrSHP+ZD
b60BIBBJCHsNr/vyA5UQ+Ojj20aKyF0cnjHqDsClqZyDoFTvJQd08wvWRvf9I4b2alYfe0FIgZnX
KYteufqSnHMKYqIN1VM+nLhtVeSBaSk/rIUFtG/tljD0mH9dLPYL8vmkmZnKYWhKJvrjH5V8FkPy
XMMG5+oQH9uiFxXKmtN/ko4K8KIDGadB+vnySzJx+JUZJlYs6XtptGHvC2M+cIvsgWx6iKZxiWDO
KuxB8T5PDiLpT7vzfmKxuG1bU2mMHpKWRBKsBa/wTtP0w+tX0310c/Tojy4wgJLQDfUQNBGmaKys
gFzOSznnklepU3yTJ4bI52hSbd8MgD4P1d0QQGGe9aLjk5WjEDY/vrqehhH8x5BgTc122PenXfZR
a7mlSzZmJEaGKvOb8nTM0wpfSkjefGkqjy3ofj/Q0alf4pt+CpC75zBnK+Ysy3XWo+i6PjtSerwb
slLTYn0G9429vt+x42SSPZoBdKNGWznMAJi8u2YL7QrEcQvC3guNn/gAjN/dkbS40EHYDDGOUWZQ
wmmP+j5V09osQLIw3EZt01hwSzSUYRFDsXv97KIvxcnzST046YED4WgIYBeJL4L5Qgby5Rvi13Ll
Bcok3l4yuLkRUSIXi/pmpivX8JalA0zWjaAjgALeHXCw58wzk8y1EpnoMrirOIPcqZVpP9CXEDby
etFpz/UXchcRlyQDSLwwc6c35qfSHbdr9axrjyvH0HfY8Kyx+3cZn2QGRyK5SrJJyi5Ch/9N3hT2
FtDT22+9Gz5Vw/8Wtd2B354X2TLmX9Ko0mMEE4o3LpPcSiqJYiIefTGShzWY4ZciICny5c55WJy/
5KREKb6u6MMNtLWbD4prDPMSQCE6/sxY1L1j6XEUaNhA5A7JNavpxCgP2W1DKPZwoA8dpmxesZTB
4IWhTY1o+2qoCT7ZA4/HF2hnQNehxnPQFLsqW83xg8DNmu4TQ4r/+pnGRsNT/glqiiseA0tba0Ne
mYdcp4Y82xLGNO/Enx5rlSTyTy/yUiXWIhLTT2voUuISLIWP8/ZQqIqxxGYL9qyQz4s/xtWrLUH3
op5y1miC2rduCmOEcLDDaHt2auh4yRjAbmVZey2ByrOunoDXdlUBierLv5vm3J9lInymXLBSv4kh
kFaTKMW4v9twoiZFYYl2AQ1oSfePucsYeDMWLFszDaYYDUv5Kg3bfCnOkN1h9IA+OkyNhJF2B1zU
3CKU0heXAEGjMD2iSE0kVEXT4ApNe2fJTe+nDBl9ili50uVFm/haLQpMNZV3wyCsVZD+l0xrxTCy
xzrxZX/UiPYII/48Q7vx07zjhrcxNOiFCJcNhYDTupua5uTlb8koECx4H45AJ1C1fIIEjsq49ss+
i+HcC6gYMv0QoM9W7MIobdo+hCVMrI4qRRZLPiviv20LIDwQ7eEYfaXCaib5zREb6bqOUU250n7W
n+N69y1RqxsHu1YlFSvYG2lwpcv3I80Ve3I4DAQ7MvBL7xbNdrXYLdZImEl0zG20xvH0pMUj0ON1
SDPdzuSXG8nHBJyidEZH5tDtTCv9NMc+e5mrKavf8eT5AG06k7CsbJPfJnQh3o3U/R4yyfyaWit9
sb5eR9rlzkOuk/AmfXAmXMc4EwxbvfLyDSgYPXVzbrSS5Pt9Dv7IOiGC8FqCEEdyvK1NVkNQgr4j
tuXP/Mh4MyqCNKDWMQUQSBK8PqBBbDYCPn1Hzlmfivl7RZRmaS+T4WdQL5ikHyKMtJXhWfqe0Y8A
KTxWIUEf/hFlFvZaWJT6Cx7I8CA2MD0thG2nW41tkFu+HOBva30rLRk0XJzHn8K0A9LtNXXIcuFK
T+1v8PDcaHxc/dhfwTwnYSB67/AIJ7hu+Axr0Mc3giMdCHwyGwt+YS0RrO1Ny8wKsR6q3auwFJxe
+jI21nt2F7O35iGrSxi4g8rIOATG9Pt2TRVybfpn+pMMFJsm8Z5T4Jwh90PcmoaaabpfjrfJTIM7
KVeHxJz2Y6VLqE+PsgyNy9ZoBqAgFlAwQqePuolmLM0RaMSlHTZV+4NTyf/w4j1LjIB/XveAndBe
Yorv9VoHvdH/9ZscFwMt1j5/EHSQzHxHX2/TMiN4oWlVT2xAlIp3gyKsatlTVaaQHT0TE40piBj6
R42VI6aiLqxgRywo091SunLvGghOTWAwE+fQ5jY/vLezaDoZno2543r2/hxulL8udH7mxjBEtLLr
FvA5imVupvG34hedNgFQG4gZIyHcchtfk7b8pGftSvmCqCNpE+zqiy2k/6xPSiKUEmJ11InsNo1s
u92BJwJsYLc2IqmyahrKfgTpa5ksTs9rcaxbF+avCpcbOOag1WYjPqPhF4e0rP3EtUlx9EvfvPrZ
njzC4oYbjnI5DisloYvsSz4jWw0i8G5SmJ5plQCjcaG94L9pGJNomPHFVdN1h1Ufz/G2fr+FcrOM
DfAxXc7ehR0+GPLKiDNNFZuvFto5QYti79gePDleJ27MYSt1B9rWVJUm6uFFwV4VNJI1C0b0IPUj
9c0OdmQa9lAwF4jBLZQ2rd2yRQFEsm4BmfbrBXH6UOS/RK3i1qKpo3hRDt6kbFxHOrKxLYFKob4p
UCtr6iiWTfydhbTuxLob3PXYpdKHLz/NbEEByb4sIJuATQ3orhzHJA0xrHspnuIC+BFcv0CQjCch
UQwfuPqNB1904r3NbhaB3PB6+rgW2RNLZwvvUAW4jp8oMaNs3cGN00Azo10oUdfil3vD7GjHRwMX
sq3Tni72Lfk/fX2CCzkCbTPcmC9Gy05B4V4n1zFSiuwtuNbRRRHesK+HdLJOuOvp+R3Yjo9lgaeh
EaKfwcA23ZDTiwbZGSCHNMiO6baZQ9NWhFfm1l/KwHKhi2GhCTqwt6z/tKBZiVKkDFt7DjWPMCet
JaK2Ore7LrQxjaoUIuHHtWPqLCq+rV5jhQd/ZIrayH93ICImgLPU76lktlor/pZfpoEsLqyLcZ6j
51Go9UdGgHMFzGSCf7gHzB+ga1HUBGheStRB3PfblA5sWQNHC4dE7dnhelEsSdsCD011G/rtWYQs
mWSJ62IdbDtIlLPg356ujzpEFVqMg9IvrGvxtPfmjbzzphXwHb7hB4c4W2fxRJ+NZXkvQIWon4cC
xQC5hVGVZIzSVHhJN0L2McvOQ2BBr78T1r6iZ+IwB+o4ysL6GDaRcgpIWqBIkm/EK6Sg5JOnXjbx
T7AdWDJns194UySYBoWkdF80Lns8xLmAJYkbbg8qmRrbu4SJrnPujqY1RvDVYNljzehfKriwwhYi
TmrslZ1uTY/u7mjbxyn/+dG5DFbaeTS8H8acQBbFuGhvokiVcRLOcMvGFldJdtjpVwmcyYA0gWMa
GnF3ND6ITL0zEwOTodgrI7OVP+arikTl3/HAtRUmiQPErN9rjwaszHwh2Key0eiq3wTZRATXC8ia
MELxNpph4hvLsqBqZf/CijTsm7ncP16LbSZotc0j0OOfAN+wxd8OG0NKBzUizVpsGT112PXZufk3
Xv6Od5ixa8Hr5t7S0EK69MU68TQ2UiXS82vVlQBg4lcn0CPdgBhtjs/fMSLXgOU25yyX4TtZgbCJ
QuHQ9B+VpPZ/miWIhs0SzVLY4ACj+5Rzazpr/IyaIn2GDvCsB/xyEIQCZPCL+w0UvZuOEJXFy4Gt
GF2fxuAYWzucwR1Il160NyIYIzVFt2S4r+S6tXpjjmissh5jqUVOGliM8vRDwj6w75Zr4s3Jmyq8
Az49tF0yq0iuSJqoKuW/k3M41obHCsLBI2MHY7io+N2DNQqVyQVqqr64/Ppa91Hxk1aUja8h/6UA
+Pkaohz7O8L/SS/X65oH7tuZ7LWEE5CVcOCDm9yeeRaJCBr5EZq0QGhagErz+jQ9nWrzBEuSRw/a
+fJVOGQmeU2Iv2NHPjrau9VFv4a8p1pZOk9CCBpgQNfhS1SceU86RtF5RIWEFQEABZvMfnKn9EsQ
OiPe66xtvi3Rk4IeqAI3fJUpZ2zot69AvP8xvX259MhVdHkaFe21bjhSEWrADyIgIhdPmMu4AA3x
kNbp15X6XiWi7gCBFO83TZL6kr2tPgrlkAnJC7Fnk2xZS7nbooqhzjMtVd3284ByVdpIsNa1fnqn
5x8xQfpDoVNWyJMn9pa9WzxGf0Ea3mrO2D9RTfrj/kWT5TnKIw1+/EhtEIj7xYmMM4Ehj+17Cj8t
iOCkYaPf4U+6C9HyKkSX7Uge4pwewfG6258q7en9dJ087Y7bLEiEwWkSPbfWyM8pJPxGO/Fn0Aqb
l/sKRYi3N+BH8IID9KZp7rnE2QYiB6C2bMTgm3ygRP5IxF+4jBrL65LVwPAV0/MIxo68DTi1jnDv
5ZhCH1uuKbP1DxX2OCmab6tBiBGScDW92JUeyXM3PbIgtKmo0oCrCr7QMfO/W3oUn/0cJEmQjpaL
DjlU32dD4DTjPaAmyVcG53xG5GBk2tXPERA4K583yiq8THQ0iSp2PbvCAzcE9BV24dmJm0vMjIiK
SWKBefTdtN5QxkbQ8EmYaelzDdxVeUqZGBEDMWQz6QBmaQB30WBLH88qD4MvxLSSfiswHnzCHvlk
LbHAIQZW0LzMBtDqVfYXYCP2qbr/5Fwwv8cmAMwoQKM5HEBslM9HLqJ+2s7mSf19d3GMzIt7SfY3
K/Q0M+AyhU9fJDeNWQX2Uc8j3CgPnL2cFdJ1U5HDRR9S9h5HCx52WQIxK+YbcpboihUiYqoXn12S
AsP9nkaicU9SS8H67DBz0asCWsU39Od102vtFbjKXur1WZJHdeipVql3grSiyn1DqiNt0UKWUcPX
Px5wn3e9aKqo3ao62PySp7FV/WguywOJzBstTFvuRdt/4TvPYPo9Ie5hQVzurvt0Z7bFQH9mEq5y
k+5+XFFbzuHRfZiwYqc4Vc8QKa/Dm0J9rj0BWeB6HYYvPPBv9rg7JDdCR9iA+vNucq9tCX0ZcIay
bPwiqbvTJYp0xbWGS6+E73xVarDAulkppsmMOMlbuRhu7ryspjbi3bnvn6MS+7+s2c7AyBI2u4rm
FiVRSR8WzVNTGRRr8glWn6FrAnRmnDNDRAoAwKmSarLD/T6CYKNYzycy3F8VgiqX1Iv5AKscFlyB
vAHweYa5rzHoqLA4eOfqzvlMyrMduw8e0vCF6I6DZ/+Hrny+Pb4K+HpLtS/5UslgMyYlBWWc6p5L
ooyaHNrBQ3UspEcmRwcXJRbbEI10TqzH8uST8o1N0QZW1n0nAz2ItnHryhFoYju4o1G7vYhWg2CZ
XC/wBlpIP6hMCmOpC4zE2BySE/hOCVmUwjkahdDaMZ2MW1NiYr/HHLFwgaugm1GMjqBiJx21S1GE
Tpwt7JR+Ws69tZ293/ET1QnfdKP2lTjyOk48pZDhutuzf/DQe/lLY70jg0hf3jfmCXlNe9VaZ6cA
t1yD4vIveg/4laTpApDR/Sy6RnEDPfBprRaicANomXu5CgrsJY83jx6VjjpX1aOaH0clxTsTDQt8
ioJCkRRXq3/RE9Uy36MlqlMj4gM0X0bPW+vrETbuK5LD93VUPPgZWBS/TR2txE/4TWAqF4qmbTxa
D4F1Uvxz9ZZxp4e7iS8b9zwqXgbKlbEn7ToCjZS/V+qmEBlhgiNZLwnP8KS7n2wIjv+TpuGWR7a3
At2BTFFjLIeIf24ymPhcBDzYwRCDS4dQ78az3aSKgy2z39kXhW5vAEdZSldN4tQmw/BFfA9tokAt
N9SdD1XJaiy5J2rxQHzv+T4xaqhcS4q/TkwzrRGY/jRoGgkvWX0w1ApKfWEqKVohBfv7+jybd+m2
iy6x0PeNdKXQWESEDu0OPIfJcq3D5kGDEne8GT4s9I0XJ1s2fKGGner0tO2q/P7U+WevhnUrTkJC
Cjag0r6OUc/zMCt/9UDe9d3th8IcL8+EGBiuo1OTMMRYsuS/JtZ/o9E+5JHfxrNaXsXVTeGBvsAp
myGhxs4OZ44PoKXvu453fiG7Xjyql6n8t1njDKV7LzYq8F1tgP4nZ8OsJ66ZMlGUNy0DIdlXwMNs
1RcDe6t6uwRjAYIUdyKWbfynZ/VyXoIoJYoUpwFD4EeWZgYgZvk+7kOskOVrgwb+5Hm+dm1h99Oe
VTUMYOzzMdPeg42wsgQrapoegyVk3eG9Iys/+Epf9kYbV3EtvgwV5weTL7DakPaWzXnZKQvIEyMt
cAAExUMzYqtJulC2+XRJi4XWwCstwTl+VogD2zjzCdj1574zcya/MgBMqvLRc4EcQnmwd3P1nQOn
jVZWf+K8yyC60a5D9jIQbK4aE1LTKKGj0NWqcVRuRRjApUB4swJttobt9T2J1nblK2iw5ekGseOl
V1hNjWLY62RmjpjbI/bYFdcme8aUBy/OUN51TDepoXSId28LZnJWxOSuEXXQLx4ua9xovlH4xyhB
ubXaJdQbr6HZd0nvHimp2Sz0+izV95lU7bI8tFpnfLlNbBXcjJ5Dhka6VGswhFZx7NbnIQTeOg6E
9p8bNY5Tcaezbb5jcY/uvJoHn4o4xKv6POsOWqXAYWFtQGnsRFlvnzx68aLzO19eJ99X42rqb3K5
zN83DT5sBaYX0/PDCFSV3ptSi01x0SbCaummP6sXU3yEod0O6ZIAGq1AaScwDDMua/kAle1otMrn
HgR3qwVPu6FrsXMDnVZLnWrDx84qZj0JNETUdpaokg6mO5eL9znowVT169P1RPNxro5fLA+c87bq
nEHFDxNknV55OmnBpPVOYrRBLBglqaIiVccYlJNWxKRaxZqZkfDPT1u41wxyVkZoHNk4BpKrriAb
xwRkAs90uRnoL2HAuE6vN7rLgMNU6emmyT8OXHGeylDEjMtsLL4I67jtwafEKRPyi+zIAk8BoErt
9J/sSPFbnq8CMclzxUuP/cd3GHszy9oZa96iqatJSUVoINORgLAGuPXLCsj/qX1qNffdCqZkrrG9
NqRuZM6iIOdD+IRQLP8iHPkLEojtfr7g7vYG3glcyQLJ1pCshkHWRhQXmpPfW3owJEwVtM2Pu5hs
YV4IuMFHqil0eUZZoPpYSTa4KC2eg5LI6RF6NXBeZcfgCKwXN97XKZDi6d2/yAyPh5tDgZJnXAB8
PFHKMLxKC4bm9vo1e7wQ8K8sYgDdnXnDPF6ompEL4ik9I6OVg5zOJ3X6z7735UJ5h2P1d+nqPnS2
d89OtNO0ClchNcF3G1S0myzRqO/lA23VUnSgWDDqoB7f20hWStuK9fnsxab51o4ZOs4D5KzKSBJ6
Dk6Bj0IjW2Ve4M/r7b1+Gh2BGrxE+2bhSV9X5gWlYtC92MgT5sr0BiOZiVtJSI40D2RA09sxqZ1B
kVaO+gZZHNXLQMIlIs6+48dH7F4lBjRNdrLwo6J6NFMBR9VpD1Qf1Ovx0PCz6XX7OLDSFMA4b/SJ
FqvGQDxFw4S2eaH23rSM5RfhYqjc8t/4heGZe9GgT+s5dK0liobDYOZsmmhODljsTeWuql7AkPbO
mkVf2DMeSFbfDepK6CF19YpsqltbplSzct4R1rXgrATvYMLzXZRYX5TrMeGvGCu8X2M4fk9a3iQ3
gvV/2uy8jLSXE6P9sgfSq2KGjacjTzBwJwV3z0+urEo3jFAVVqHi8kVxqYx7lXd4C0Eox6wFqAzX
hJbQinE7gMD8L6AjCTxj825veA1aXvHsWyXrrp11IRakYlbalxRlVc/SkkXKIxQeDgYZxg90ggHV
/eNpeu2KlNkoZbwWzltG4kzt294Kg6oSJJpjibrSeUqnJeyIJ9xOMNk5jBMdvj/3oue3QO2Yeycp
vnAeqcrplMFy3OSzx2GQh8VKK3Fw6Crzny1XRyhdg8qehjaX2uVcrsZwO7/dwY9sKJlpw+dYqeue
wMwSnuVnO88LKRpzOhJeXEZzEncyKD0P1XzKGDnRpBXwv+UZe5/aYrBH+sk4VU2YuCrV5i6Mmw45
of8L7rZBNDjfg/1pBZp+r25W2Qw6SxrMEUOM89tKusTqw5bvnL1Wf29mbLeU1NVtBez0dtZdiOB0
Ko1QfF3AqDZG/Oe8jCKe1+ZSD1GJdP3XvdmUlpohun1JcoOnuRz9N6BsdAjMwPU8DNAyyZxr6uvW
4mB5YU2MhnM2GQzCmvKznpqlPm3+ypRH2tUMD20XByIXMSIyz8w4PNBWJMn+wXgv60RHcE9tKODE
2JcThyIJPcXPKzbof4xs2adk0ifR5+0vJZ9KJQqWoyldhLCstq5tJVOy1ig3vpvKPHo8aQuPcsA2
pp4yBxShHdgi8RUX4pH1CRLzlB1k3m8B72qGyYxboU6H3E4t4LCI6XyuczlOwGA0GxPzEYX0QDgl
RngpF4JAnLJxalIPOu8KoC/2tj/nI3hmpjBSw6ID1oMH19jwYUThWTa13K948wP9VcbpMWkvZWHn
uUNVWxCkB8Qbg0aH06H44D+73DmsYiEILlwXUk9kZEXzlMt8EyUD7ZGzOHHGI6k6YFdu/a/zNXni
CbgvKJ8QLZyQgbx0tj7a5+eAKhmiJguKA1GyqjBf+r/QNj+zTNXK3+zXgYMBwbv1qUXhrScK++2B
rc8RDA/atJKg+LfFoJfcJWuAFK8xNiN7imehZDaZ2P3K+8aKn5mGB8V09EVeqvRDyGlVIVD0/YQQ
9lruI/OfYtY5PiXxFoKtRcJm2s7hVCn68aBNxbLrzwA1fPG2aM3fqi4B+AOggk54vsLaq3ShHEcp
E+piH2wD8xXClXpZq/AVmTl5bb+mZEpkpxWJJpZaYzbvEncNJ7Awx4/heoR2rCQ57sxf7ASz3hrY
koD7uDzOe3absBwLxlr3xw6PU06jNxB0PmfQg6nhedUt5KWCl8f1W8ikuF9uZrBnfT2udJ8cflB5
VTF8Tfuxn0sqkyNQFR6oTlJ2H2a3zG7CUwHuROIFEvmjlMmUEV3ZQL0Lw9IvTU0nUsIvj3dV5chV
YW1aJfVUTht9QxCiQSbFzjgZhN3oH//lGfaD7sGFkEKcnOI+sVMXrp6FvYYnHmDMht4r/Hjc8ZHK
izhdh685CGI048XR0CZ6m/yhVdNBuv+B/qPk4zPV/z0f434YAJpm+IZJSTL62Al/8tzozXIcJ8Rx
s/kjHg6c025WBz7ciW5fsbaOLi17Auj5EKf+Ws2mA9Ejg94xRiEwYswGKuGW1UOxjjUKdI8GHOZl
zuqQiAiah+2SpVEO2l2C/MVqgCUT5TXgMMcDwB2qZ66mySuR5SK7GNbjlxMv4efQS5LYsvJ8DCSp
cY2cN+6GCBFeKmPLUW4st1rt6GG2hiYYYMu5psqHAsiNi+sBwh/slDB2bsd3B8XzTGg6oT9PmErv
Zqw6liHKO/ScajRMc7IxIQlm7605cZliVfeoyB/2yMwigtmuJ4CQuBPRYle5WeJNwzVTp0x7NmRe
CVU/Sqo8i03EDX+AL9UAm6NjtCE/JPFOc7qrhh+26NTI6q7ZzrQSD/GwJdvq1oqwfsNH23CQq6Yk
NQf2ejFU0b5Hp8tNxjAweoxoELpptYkb0Q0ssZZGIbeiQtz+n2uvGifMcWvHpg80cdAmGl1d/s12
gR8W+F8B+wTMn3e67mPop9QiKRl/do3sJ4xoxyUCeKDgLzOTBJSJ65grG024gqPNp2TG4YWmYeh6
9ereu50nZEjFG6KkoLfpQCjK6XTqtr9KAafFkR5WK5AUOhoKeXz7ShXx6sTslcbxy77lNhO/cl4E
BETOclguAouruTXJtvsSCyxIQRmB57v9FAPn5q+XX4SbxTcOAy8cRW4JHF+WqHTw7nm+5Ky52QzM
M8xOB/LT7Nk8SluBe/1W6iewrpJQFcmIE6nuI06A7fS0Ce5JCEddSTlUDRXa1J0S9vz+p3KD4eAb
DgwjYU5QDo0bplkjl0JrpzK2mAmFCKvNsW8AA71/5Fpmu+a1QcSezVSKzaE4WDbn/i/ZCtWXBSB9
TdqDnESz/f+xds71LvjX4O4cUp2HmeOkJZt/qVVW0KgeNA3O5jLuyKxpyflUhBt1NdQu3yk+/aMG
18m/ibf764PzTaSA+PjxrRegdsuf0kZdOB052q6Y8I7jEiZJl11x0/rmlGnl24Zg2eyzYM0IqEXE
D1eYzu8khhM68QG1VeMyH5usqz6jjHSzn9ZYU3xdJkduxCV8HOKj06xvy4Yo4ct/dXXy//H2Fnct
8WoDNMThTVs9A21o29YBe4E4gcAH2gqm4IOVYynGl4pB3EeL1+d/2POuZvAkQDMkb8MsS/t6crQN
uv1ld/UVO/X6OxbrS76brFmNTlT92QqRzyE3knxfxCwZ1kpoDU+ZOgSVjhGxx8W0V/YgVnWPy8S+
wB53OafczUpPQW8E/mjD3hVaKyzxgr1EapIiHDGbvwRxkakWP8+jpZEODPyz5a9rum57FIz4+A2p
roVkfaw0JshE7C7WSNMaERBgofpRR4X5RpqF/ra0N9uR8Dse8P5Uvf7vE5kyBCiGJ5KKFtKH++70
pUsw9vZWeDrSnl6oQ0lCfQFe3tjxdQJrOcdlBLVMPRUzCMfXam1tU/D7Zod7xW5QqTqXRuMqy/HB
XUMdXaUZKvQ+MRqWOAdxahWjyJ5CQdIh1ekAU6QHylF0qUKwQwKMuzLcVBCFSZpkc/6aBioeCHG0
4fkQ+p4b7Rm6kyUq1AXVDnt/yODElxUEaAQ268ErsZs6UzTrteSKeTgRnybDQ+fG9JFxzqO8/xJ5
yOVtUjRqiC53djU2mDXqd8tfxJJlzRkyh7/AguEMBIY1CdV7HOrXsCE2nCVmPCKJeuY+JRgE7whL
zx4nfPjGWTwWYhiIljMbKoCjTwxe8M5j/qG391zTe69ZfF6uGsWub3XR+v62qJbYvftVOd3ChBtS
p6d9hwiepTFsNlHWZBo1DEki0321XGlCHyIlyQXJRxANRBQpFNx/ssoc21FVk/9YNskZzL7sQrqk
i+fFqw3Vquldy5Sblf4C2aPdt3xeDXchoF+NQPiax5Ty/IBY1XCDKWVli2/Fp1qS2e43unF6dHfe
p8bTyQo4j/5u4cSEPyEYAQlWxKTsnrJKky6wl9qayXpcj3oFx/amzB4KfyqoITyAXuwmyHfwgNUe
AzVWse5mGpq/bV4uDeD02R2qx2E7MDuaX+d4sEiI1Ygg6cGWj/x5h0MZ4u0bajUi4+cZlT1xjlkt
Lrmg+sEIadfIP+ej8kQX/LeBza5lGQaVg5ydsV0WniFTQtHUD+JhLoHBIZmX9ZGlPedlED9bfIiH
GAaN6Hur0JQc+F1XtoYYba2XV5HujL6PwKtClRa0aQ7RTo3fbxw3ZUoKlUGh4YZh+vvCSYjZ45Hl
ZXMEtOvcqdxE45+EkdnXt4boxzzKsmJMnZVVWECew6UpOLWRma/wKHxmF4N2wA0ktfV89EALum5o
OxbWrlvu+Q4PFuHEwGV8gNBm6qVomS6q17plwXRUgWPQNKvlWqiF9puZZ+ZvMEJVdIxOIqlCFDnc
vKYmKiwFDGkHc+lJewhFMdyUDdksQFLKpFlcul4bm/ruHbkKCnVqN1OnvjHkCiCOV3hayIWHlbh9
xGbU7p05rf8ctkcKmowsgKNMM2zHItYVMcJYCvhjjU1x/zN0raNcmI/f4FDqs96SHcpkZRgzMiGu
F6nZ4JWAuTjt26GELV/DJZWavmpG36bXkIPN2sBOkz8ETCug5aEP86T73QHLgghgrZyGNGN+oTTY
VfY3++ymMe86KoeYu5k18R2L7obAcwd22riyWT7nfywgU1li4MDqLUT7fFusikY1vKQYpqNmY5Dg
083aj9hzgPAUVX/qTRtSMG/JJrkO8j1YPpZV4xU3EdJK93JxtkTPq+7S1A9DMql6QncYoy+UI98a
wSZnKRtetETm/OW/UTL7U870Ge0UKvb+7XRrllxynGTa5VEmGOFVyLxeI1oIukrFwJ+hulEplY8k
qJjjJuAcKgvuUavcU8TbOYZGCqeM2Uck4B9+J7LDBOpEg2k1fRnDMfiFTLnzhygI3Ziz5B/WR2Jx
bV1xe2qa4zwakNHAsTD0B8jLkG97cE6cekfkdrZymFD/bTUdd0JumkkRmFbwv6WxcWOB/mvPNcbA
5r+s21Qveg+QaYU63fclWk7cnum4rrfduSwuX/afCzrAq51DjOLVQqvijo+bd7v+tZP+uDYEeIs9
TXPGEnIXf8o811ywHSwsRhb6ZuhHg2+nO7y+fCK5SpddUnx1YMl41vLilQJsZbiUyBZw6JbNqT3p
eJVV905x1AWQ4xIokPndj1VOJh7Vb+iy5br/26fGQW5qJGjndX9DeXCSwZtJuLIG2Fkyf3DAMNp0
LpD8vcXP77DTpHLq+y4e+GxWs21MhusOBGguBM95+Jr9Rg2DwI0nwNu8TUkRsMw9YvgPdB2AczGX
ZR69+MKecy4YbL3GgQXjvu7uibTr9/QHjyq1ZH63+9zUGwoTCv3V6oFultkStOsJpRWNZHDnhqOp
puqYlhXyhJL/uXIwz9i70zTltwahvZj/o/64SLZKP6FwbVh0zNSQNdoGrz9nLysngCnsBwBS2z9D
6FKkf9qkSaVEo7KG4+zRbmyHqMV86IpRXat6xbwk1sQljmoc69XlD8xGF86gddwTVSuVGFeemOG5
PRvHfaGI0Co3Z43WmpqOG86LvQrAeFyHS49enzvd4Uv/VZs372qdmHllVHKhX1VRjd784LvmTspY
uIAv3GAyWrAVLcnLxSVJJUD46klHFQV5X9/FW9RkT06DDZBmEwYejxkJ8k8EUkYo46GIku1hLXYF
YFYIwJ3fb8vK2qibAf6KRxoWbPrE67RErngGh3oiLYv0X0wiDSh+gqvVXAWr7+X9maFa7ZX7fLf2
OCTaiuRdsSQSV7YRe6jlUX39GsrwheKqV/ZP56e5kkN6KmjQghdbmi5NcV3qda8Vyilq4G9Owk/n
NOtJ181emcs/QqczhWp/bk1XkoJimu1U7qdYAuXj550um+PlY35IhJNIiqDRgSMmoZwQjm5dmbrs
unttJ1QoKCuQmtWUJpp8gV/I1jS5VbXE4p6odwAs02Mqs+IVz20z/YXWhGWXTydHv5LfxIByC+Su
AhgrnyxTV4qLx07hF6Sh9jJCwFdfEe6zAoRJ1J3cp0xyUKWlfImYljt0AoOjLuowGiRvBIjkijgk
N23CfiTw/1R4qemepX3OLpNbS2X86vUc8/yg6JqLEZR3SP+1HJ8EXY1Y5Ze8W4JaCk+S54PZswbF
872JvQjm1r+9ZGncWxo7/LXIRd0jQEmq9w0NPG72hdeLsQmjd/wR5skh5cEsp3G25HswU6bdAf0y
nxP9LIhK9w81h2i+zLOlShsu4vkVHVo0csF8kl6f0mxZLIm8d7+hyksW6Lgwa1JJJqQw4Fn6eOSD
mv0PhzV2QieYjoBK9ZGQfdd0/OmIGxPJlH62gDDJAz57kvbzudCkfdB/dYIc8lYsjN42J0hUWzKf
2xNYqUv9123I9skBkfZl66Pb4CDn//gLQmNTxdALj3q92OkEJJY3Mct1E/DH7ojJ/r2xpWwirI81
nQcTRBcCffhQJX1UTJQrC8nq3LDW90V5pUCOrGz4V2X5cOximyJx+65Jx6Vk+m989xwpCIe4kKst
098MV7EuW+9Ytq/zJek6zoAvdA4ReAj664TL7h/sz7hj4riuhfsV8tqcPfAGAHScwg+4ere9/7j+
dQL7+2DfRrTTTu9bg8ej6pXOIN/Ny3+ys/kjZhcEu56GqQ2z1a8IKr/4FMVLSU4BpN6CkqaK6vno
Il+Xq4CPytGvV/zTldJ0VMTRR6/wnXOFhi5pXt1Pi2Z1G5V5m1XAJPzflTO0Qz4gXiQSLbOPNyRY
P5wo1hMYeJiNZ2Ha0zpNHGh9TSbpy0T/1GZ1EqaGvb6KRxCzULUv7YpL7q6FbnwkekYp9P8/xyZg
A1TSsR9XABY0d48Ev2wIOvwrcifH1pH32dGntrRgYDYx6NEEYBTbd4lXcqRl23L/G8NE8tfysGUn
MROHPB1H9tjJiV1EuOoFkLfooWIdBdsXklXyQyZvtvKObxfyoQG31N9t0FX+YZO85cJO1KXhO2P9
AQykndvQWVLNeCskBA/3BHwGCyGij40TYB8Z9cRUpYUpIwclji/qrq/3UJi54mlMB37zg4huzdfY
NDC3fK9uDyKm4c7BHi4zQaMDiG1DnQrmsp6quctu9PM5ScUbZp3+A9ni7su+efMatZ49r+qtazIa
A6v0hDg4x2Mv5cxeM5oiolAzFNdYzRljDw0rJYN3jSwtquOKR5zA2/ARwFQT7wVng6ZR9Pon7BBa
NlzlbVexwyqOCdzDmpexuqFyB8eGFdJ0UmBKCjwah2Nm0B918TPH9fW9gg1tGFX61TqDUO6qrbvw
0IfK2Osy5ARPKmrBq3FFHcEAT9eebx/2FSP6ljc8jsqDAXXFI0dtOcZ3LThPyc37m+/yCOr7cgw/
2jWwcqQu6JoBIKF8qKWSS/3IGfKPMDEv18Jk0lVH4ilOsUO5vYT8IBYqJZ6bQOEkt7aMDQD42G3q
Vqdnu1aa6qr98KBFheBkkLcffDlu/mePBEuXVWz5VEHLMX42hVjsYwzrAQLl6RLzV/hTvHngw8+F
TvccKy71Ssqd6z/+f65a9+3kVgM8E2iZHom9WnESflia5rPhD1WjIXJhrPgrFvYZJfQuf1N8TklT
asOOloQ5BTiivUhq1h0oSzqnRskTmVSv8Q5dNcOFQuZL4IscL9Kl0TlIvV6V2Q1B6mV2oZ7XtcRF
W2tHhUQYBFfzUQ3cdF77n4oZ29oq8/9YdiTPPQAvXkf6qytNBLnR2UnniJa6DYspXBm+nVVCk0WE
IruLTGKKWL0SLionUanQTNWhLgRm48hWAkjIQyhCigzL3coo3ujUhSXzoMHkhpwcj5t2bxSNvFLn
KB21EWoHHa4FIDj97l0jd7AOtMhz8l7phIevDMWDh0Ty65UFFNlz08OE0Le3NgvbRk/q8lgnmegi
uvoFbACWGm0WLGtgGaHqevzY6A4UEyT52tT0XH0kem/DXPxMId51NGpqM8wR6EHMzTZ4jJCO60ZV
voPqF+yYe3/WcGTjISKA4I9iTyAAsCa7y39t4ThF2nwZqZlj0ghlO3R+BW9+1xKeml/lcIk+K8dk
bEB1H3hXvSG/eyPwKqESO8UMY10nLemFoEFMXB284ZtJhfvhmQ40U0SgxG7J/vIxoslR/vwl8Ym5
n8FtrzZ3UqBz078WGR5egCzobd7S87IwvopqPQUDnLWWPWZ2hwr8Gwvdk82vwvCVmAl3pN3D93Dt
c42NKbJ2uc0Pd+siBWxB7EFwQQMWagLdLGJEAmQTzTQbCh6ajMDgFWJofdAroJ9yTeKXmB6zBFfL
Rp9veZmTFTMFkiLSxVqqtsWzC8BJs14RmEm9H41jyB0hMU++VmvKTplr00zslxQz5nrF4kquwOBT
RVagJekBvadQyIZPmFqd1rUf84kksbYkEchhY0J6d8eniT3ACrksWhgTUIzpckh9Kw5FCZCVYGMh
eqX3M53sDDdbAxog+Ed/OZr9kqCKZIKJUmh2bSKtQ3XtJCyiwzg8nkf1LnfGthBnOYnTg3hDqa9I
mBbL4ZNthGhiMoCL2AlkmmuZEuSsyI6wD3ICNd5PLDgPsN0v1iE2gvxRe0dA0pcS8Xm02ssjUO2N
aN3xIDVmpVWu1esuvqSwBFaXMx32NAfNYqnIZVsGJEFlbgfbKGKrrvhN0+2Vqb0aPW62i/neTilL
kMqF5YGTY6d5cCvyBa7mYcMnF6U1TgEA6WgNmiXGopZ//BPpfED5qIijFzkuBHXZNGTYl93AM9xe
qSJ60YtmAL6pigWe/6s79uOYprb0iFVrynktKH4NBkKYbgefnjdjfoWAIdT+KbhIGQ3MuC27a+n0
/SM5+qj6bZyx6n7mMMGPCVj41FWCTnJefj3GtB76IHei9mLwhRfanxAYLhDexdjY/cSW9/DB4Fx4
UH5GGSHK3O35qtuI2qrGCWR6wLxzRa+f/QwC3qBDy2XmbEB0o0jP/pdNAdPKfeNe8cmN6mLQ12Ms
XK9IM8tTdxx7+FDv6pJrJlEHxfVb27PPOwXRy/UPQrRJDipM05EnMk27XXpO045T/lxKpdquKB0f
npOgNtj/5u8B0Mnn6YKjiavb68tNkLjC1bdyOjK7noiJreBn4fkuEBf+aVBolQwWd+jY8tZCH7cT
zo4Z4dcRv1pIzrcflUW+kodrQ1+og3Mh4/24hcvMAeCHLJk+uIoaBIU0++xBiwQXwy+2ySb0t97D
HsgfneRUWpoAqYmv88g9+8DrfDT9KvnbJLabEZygAShzeAVD4TTmQ69Ri9R0zKrNvAzk7z1ZluSI
hqM3p+aPyf8KSbdNZz+1DkaA8veepQy3f3f3br+VxtWJE45yl/ptvK+b7DZMsUkxYGOJ3+pssC/k
ap+SSCwY7Zw6fHilPpoUPcKzSb+hyXFecbWdv4XIRBWZbjraWapdBA5MfOHK+S13OV5qxDMoeBfK
th4ROcSdh8mwoyAG9zQ71iqGqtJ3OjgIngebpMkO+R+ci/Y2c7i37FXLsbgGaNRGotVNt3hlrtLV
ca5ktApkPQFQeqXS/ECkS/PDb87eSJyiy7n8N0fA/n4ViSHcdbjse5fKJA4Yv/TY1SaUPudsFEgS
dfi20LL49wbNTxk0tFL5wK6jp8bk0vyBoZ5f1iXHBdUOnSdXtNtd1I0+do6pYnu6+BalyNTnYRa3
8DFmCq+aYy8TOR1RKkUGBsQbJkVxaCTxSNGtIu3WXSZETWxqNszSYNG0Rp3d8gq6ybvBLHyRdEJE
jh8XrbScxkuKPkUedaWugr9O6OgakaM8bSjoVI8yL827Hd771GImkyS7b9AfZsngZSHUN6KejmkC
6iFr/b+A68xxs7zxXvWN4PlY7riALPBOZzMpsIUk09UOWkcZbLDE2nmHvmCijjoVPebO9NHkAsyT
ozOpM5TArjegJOROL7d9nMrf7dRSjH22Rr0qI4YAkK/mJP9lt2MrjSjE5++quX1GqSsvx8/jT0Of
jTcLkOsVkvWb1LzFDyyBfPSiUG3+uFLaPwWG7YxPwIahIMPKln4Gkeoq5fsgdfCVpjxvsXS9hQ0O
hRwbGOqxgdL4DzdErHi6hCoLB938YBhnyPKjw0haZ+CeSXfxOrZ0SLCFzqxfsn3JLE12PifjdujQ
YzVBevf9w8ayWb30L4ARIHXljqwTxKfQa2JKzwQkQqyTAWUNVcYc/xdemmJzFQ7o5Zchwvf01FnP
XJBd5jiHk8MRFOQFBF1CD9RvwfDWupatndPr31/2DGo+FcYpESqyh8PusSpOu2kUN1x4bA2/w8Su
q4KhqEjUHqeNDPXR5d3GOIimd9SbzXJYrtTvfzeD7hPnjUjMofAMPz5HmtZn0BQ6v5cojPa/jL9q
7xBmf793bSdDyQZwRzT1rTYKuM0XHtwwe9YHLLJeFxnMJcytU9xYjK22oRhJK2LhcD8Kfiofiqip
kuVImtkcylR6UaHzx5SPyN4AEtIJWIv8nAfim4MiUCH2E7DQiUwfzp64qvqXxSJT+RwRWsoiDMjj
xcOwZWJAQTfGFDUxvlJgbCLVmQKyiiNg4ftLxC/CPwnBAB1HMb5vsphXAor8LA25GUV1qv8yKlFj
PzgfYPQqr/86Uu1MyKoUy8dQA32swjoyBg9s6bbkW5zEV0COukamfcoS+n9NEFpaUXE9P7qCrUf1
lFQE4OFGfHRJ6B7UiM1NBU2UJAlrYxGI3d+Mj8FKE5oDhkJvT1WhaHGmtNOSD9R3ENi8YmVR3Pf0
AyGTzIrXfnwa7F7EEhEleCdpG9x41b62y7dNiPnoxmRLURMgklwV3aN9fHLtrLMHeqD1vx4h2m7/
V9hFeLHgcmKNx4lCyTy4FV29Tcosno8WJviI80ysDPLWknmFWBJl2bFUd+6/12tcjFsQzmPcERt8
9l4dqxuf8J0hjR0Y3B3QXs/rRnEtxWn47TrNHBVSq1HM1Xl/O12a+1eIfnZjdWa+U1/lyGm+W5uX
+DIzEh0x6aq0G2BlqZMv68H4edOLv6XTAB/2Idm0HoDvgYl0lRgFOoteVCAX8sUyfR0gdg/bWTOd
fjPUxrhg/7BxWvOgm3xdiFZo3OPTYAOxHqzgaoZwKgwppStgjTJhyfP+ZPDw1TpT5s7v3d4buCv8
XrSAw9zbL398nXu7MC0nbrosw7dUDLTEywaYWxIuhbgj5B3hPvpl0l4tjQB5IZ/RbGuc+NbA7stR
sEeEfB5yERwKu2EFWtJff+PCYAr3vnV3dWu0lFmuFLbBgwk7CG3sMAiuLvar9aweyey+fhteRZPx
9aGCmzXSsloolOKlqWE6VPbfiq3WoSXXi/4g/IDo6ecSm6VO//Wx/H5THkKJyKrVvMFHcE5dIZvT
gc+GXPsfiWRc0qnXmrqbAWULhwiqrby1NcvOuQYe5LV1knm2/rpTTiTnlfcaOx7TxhAgQS5qJUnX
VYE3n3oRo2/eOvfNV7kJ5GYkDNStGY0EutHF8yNM2FuEqo1DVciU06P+F1Zsn6IycTpIVaNkedGU
QeaYHDP/z1GCeWAL5qTJR8Mo7REmCayCvXUG4p0PtGdaxjqBxJURkaPkeInDZ2ivDhsRTiSrywlf
vQN2bfA+L3H2xMfQLwuup7RANWciJ4uGQZ2Udo9NAml2pbvE4P5PBDyO+Yv1TnkG1L/4xLjw+Bk+
KZ8nEAICVGQJZxzP6GHJdA+m3c2p7WY7ShpzMlD/PEUK/P9zS6blLeqZ0YPl03/v1xrfCT9IWsZb
b9qABxu/QWYywFcBkox9ccF8Pp9zJtw+A902idujsL5dQN2/UK237gxCScfFF82feHpjSUYwR3Ng
K35z55ULlMkm0DlCA8niGwpdhjRYXxi5APY/F8X4h6iplacbu68QKmKEOGklpx1cltqKKKzkBqK8
DNth6JcyswEJCmb+yJnaTqE71h6m5E8Bv2crKPc8edqk9HmKQ1EpY13JUT8R9HwkLZfN1dq/yCf4
CsFdLVhOhu58ze9k63oW+s+wqBCyI6LddMpLwXDPOUswoDPQFsGsj0flHftP6+nJ9UPXKYHDp47u
0prVI/tjXc+hjbFZPfQiItwP/R09Gt8ALthzs6wcuY3JQj+qxeXRQOcFFG5yd0Nfpx3/8XKOHRir
EH+Ha+PdA8yTGRIHYOWxivTH/ddhJ79elU97R6ztS7veDXsHkUorq83tsRo/WhMU7aYllAk85Lv4
afffJlC6/MwVEwE/1WQcx5RmPcN4jvQlqTwLDYCv/aBhS7AbqzBdhMJzkXk/O0T8J7lbAhSsjk/2
uaYLf+CdwiEsc4juEUU8DNUqvC/zpPHnj8mBOJCILkA3H7Z4U1SLyZn/MAwFUmucQ+cn1fDGO/Q8
HNkCWB/SUpmjLEFQVSL8D41TFtjZBN9IVmC4LlpLj3FqFWlwbSKsZerDNCTZHCTBYb+Og3hj4ZT3
6UD9fvdf1rrrxnfjDSnXCi7AMgiWGLcvgHMzQonA7QaUjn5mJv+NSViMB0Af3KKigtCH/GjJOJob
paiX4O5zgRhnjJaFzRdNZQ5aAx7+VAiFrLaOvOv/5cYtj+rzhtWNK2CsrR46A6q8gWoLH3AjrWsW
eK8sOaxKph1vlKq6aYi31g5tJqKyWb1phegLC87fPu5MPmtd8XMjCQ4iBIRfoTLaggkMwo+eRQHj
G5KexTBu7I3InaClFgmy100vzIcNAg2zTaj0Uobrib3OlZ94mwCTDYP6DPQJ/9d80By11igJTR4S
PiprBDdrYcQezUrSoFWpkAPb0FyICyNt2kNLN3AktRcToD0XGbyrBXE4qetKNOQuGN8alf1QSOmU
rWZWWLEyblYJvwmuIA79UKwcS04Pdlbf7umREsrvpsA7WDKND3wIKsz+rYv7ccbWhvUO/1M8HvLF
VLu7eKXRMWqES6kDNUjFYsN7sstl1MoqrqQr115bfoToB5ScFnJ5j+CMEQ0/5dHRsy1HpJ/iKqaP
Uag02Whflq6aUzPUZJkMf64cp/NyFx99rPdD0CMbbJcU4sNAKbgWvvG0eIwNOp8PMwavUjntbDLT
j3/GrsSreoN0mrGcMyp+RYJa8GpBio4Uskb0o0BWdnFZP07dOrI7CdgrZyh37qAAjYp+DL8vizzH
PFt7Me1XAJKDfHw2VdrznrIXBnsX+3+uYf5AGBj8u31OJ0e6/GNN2u2uMJI+etrZgvTHi51zwd6m
gOPBi5OimsQe1AZLSLFWdfSdHQQE2EJZUDB3XP9nU3/rxkSP64gsz3eGJp6d2wGK7D1c3xWPO5l2
4X6VyTjFEfL/N/IzCLXAkzKdoBrkjma9d0b3ZaIiH1dnfBwLsDBhRG9qtUUtplqLqFSRl8l9hqDW
ujB67t+CDMeT+E/iVCe3F+AKwiZ4FAQX+zuRO9YfT7BtTMl0AP4m4wq6nZ2y0EipDQHL7krJQnE6
wQwSRdSAr4oBmEX+YylFfVh81xVBsjxLRCBJ9ztc3QUpMW7aZnMgsz0gkKPaZ9GHGjyQlBbF5k2K
d5ScNDnvpDyzgdtSuxZq2wApLa6csIizlv7ckUwtLS6h+iMJAz3pmXyNIoLdWb01UD34Wvi95s4T
arAGhjwPTrLcyEvWW91+C7wdkNJo+Xc39X0g4DefrxN6ZiWltnMI1d0uQUwcyyCxaMqG1+f9Sjsg
ispmio8C1g/mOLOW11pGWgebl2Fc/ntkCw5wlFYM/kFU3yT5VOSxpOeUc9A4npY7ykezo49xEk3l
8MjVmJKBTX0sAfeUG1o1awzju4wFXxtBFRkBMnSF83PV04JGqUUvVtXx39aeYJ0swbDs5UTd1my+
I6SDhHcIO91k820E8kRh3vO6rQCgF5GxOqFa8jNjlnExPfILiiWF5ic4bcdlresogugf028wud9G
cCbpZufUcx6uISNZGMyYqybQ39QckWfl4w1l9e6KHXAd1p7z/0KqUJXaC/8r4J6cxFhFzrlf+lGB
A+8927F8bTYf4DRNmUIr2jdVnw+jXqXItQiruIzLDKxNvqUsv77cBIjfA6WTJQG5mJsBn/tZVfRX
P9PxJKyFGMVOetot9badbmwuVn+vmeEE3s3CSKLmRhZFszfw5qa8gUdyi9jgct+fpPRsZxDoGe7F
YOcF9AMJfLq0SJjH7XcoI4Bwgir0NK2AboIpmD+WeBOzhfEBcTPlhagmb3TXyoQ0wYwNpllqzL+v
IJiNxAtiAz7k/N4mv7pk7zletaL7mtQVw832/ZtylIPvSJnKXNDKYBHDhWMKDmFWgA9JkG9QAn/j
KyGp0yEPoLcM00QjXL2W7FMO9NiXxZyMiwKwAJzWkOw+fFStKynHFqal9f7mE+UGOZ7TZOqFGWNb
AjPcAqPR1yxN+7ntrzsPG4u6FO+iZ4gpvcD9mHPl9W7w9UDdU6ZEoNTghl8pdy8XZmakQxfR9Ujx
Z0QP8Y0KOSsiFhntr/VJ3812tIA6hj88Li8l99M3WYfEUXuGQCClX8Jnpz/AWt+nyeYR1+EPJQLx
MPRQGxXOvXKVq6SeTL+LIkLJRuomiwIOnnTpo5w7cTo6AQZjXkdGovj8mmwle9oVZ/8+qmAfW7y+
DBzUmWIPCsnecXlEjgbqNnt3p5yXiuhhbtmy49MEDggKRCOauZlK9OF1XpuII6ZQsOugZKegdMcm
dbv9QF6t9O9ZS+5gOnrjTO0NTD0olLJYYiEyXNqPdcHAKsCRvKxpSceDb974nrwMmHDaB8fE9r1H
1aWt9DAs35spT/QYzivXLhcT0wHBh0p7ZAd83MS+OPf6lAANNejqElto6fIkDd0nb4nyohYlKIlS
QgJcGcYK2hQ7Ye4kMTTCBIZiseWKBxUAYifTefSvjXPbNpKioyLTn0HIZpMt3oNAUshRzKdC+cvM
2V5M3qkTIsKDodyWOSKGxIYmO9RTNEslwDYiDhW8Nt8ImEvqc9vyt5VeTUUGK6UEShRC1KzbfRGG
45OUCMXj2CHJVKgYINNyGPbCLYmU1YrwvOmbujneh8DUkm4OBxMdA2shBY+edPA1EB3+Qvb+Zxgo
kNpT4XgusNPO/zIs+H2ZuPCZHezASpIPYgG5KMeQKzytC/1gjNvGtW+uJS5HxnwDMNb334KE1ytW
3w81xVWlhhtYtsYf4hp/9b/tHbLNkrYMHBOSosG/irAWDoQUvLI4HWeRIAIZYjUjEapm+wz7SZ3T
Xq3mkE1UJuXGqneaeNpzuWFmSMcIWZyBKt+q0YWkms3yd3DCa7RIdWmzqFya3tuXBi7LoqWvqQTG
450agnsOm+ZBtVIx2RTYaTquRaKGxWEMucNak6UNcL92IoIYWY577QkGS2cAJ6TFMId2Nfx8LqwW
0augO8XthI06rkWPwaWtcRtDolEMNNxQ2s8YJHGH5n8Mn8VHNDrfFKU4xBwutdo7SpMu8zubzBKp
ZYNDJfipmmtfRbL48xD/oaRnw2decvLP4BPyd/eo18A2OeKLOWCCtM9an8ZX0dol+p0eK8+eqHRr
sbw74bWKXu1sc+VtdfzlRgI2SZruZSw6OvX2RUo3acufdkPxPsR2/tysE8p4KJ8yBGviJMtZYFFn
i58H9L77qe5//gRHfXVv1IgVKDJ5nwzpgumipqlNfXMznW3UwAp+YuQeLGRjjiNfMTN2zvpPfam0
wX402uNRvubOYv/T6cvoSm5i1qmkVXRfjGzGS3MPWpE2ha7Muu5lZR545Ak89/OYNacTWsQB7l9A
RvLJn3ZuP1GIkLCVmr0Ug6D016B4sqnXfyXJnbdJTJv/7NHCR0eftI7A9MV0p9LFMkdah2VvSfUr
rr7cbYqf3RmziwIC9I0g8cgng01vOO+g7KAIvYxq2kJIJPhB8gB6xjqUrBGKTBnbmsZzQVp1TbdI
gCXmG5SmUYOZi63vwEg8s6R7oH/F7OasjJa0FzLvpv+Nn8AhFCLb28kh8itVGGl5mSMpb2PDqO9X
jYSjo6drKNm2TuzCqdPW+YppOtNuJDVNztQIVtnUHDoo5TtITHqaYahcnyVV2bTmFXU4/lHaiUHc
DU7bMdrVHVoGokPGN99VIxBcExjIbfT4rqsyVh9fOShLHehRDPuqtCRkS/4cS5048EBpjbMaOrQJ
bcKRG6XnbYI8RiS044eFbUMLij4lqPhUszXF3g6yw/bDFPNfJwc0W0cg5Jx8P4yxSu+BdJGqjqv3
EWog2gN5UEWScKNZFude+5s/9a4stk59C52Wo0AN8Ccf02C5QJNkUhr1VjL3b5H6d+ZD3HvUkhLj
B2QHIih6E9UV3ZOzXt3tnglTCEh13I4emyiugtYveTOzj98hS9LSGrKZeNwEMpowd1cob1qo84Gt
NZW/h+Z+HTLomoOWZ8C76EFdBKyuPcOoaDJgBAwv17kIS/s14CM8u9/1DxsKu/YOEow3Af4dtnKu
K8wVBUW74DKH9071QSyrqNgrA6z/f9eqop3morBxHC6MRdByo9gFhEgEx8vkzC38YRBxBUoOGtKR
3HV9GVFdo3JNQPG8wsE+G6u9lH3ag7ZlXVAHhTi6Mq2COjBiwQgLth5Ffn2YM4pkQdyczI/1ecx8
gJMOWlxEmjaIrYERUmrwcYgQC+/oto1OMsHREAsqQPC8Z5KmuTkLQGPS9ZjTGWwk8wB9zNxC619n
tsezF9/o5yCwgSpTRA+k1Ix9lUbvvQOUQVxDQ+iNPlaMvu+EF1w9PmRNhVgGLYhvnajGH4d00u4T
snFVEt0LWCoej0oDpvJwM4Yhlm6TQi346/pKBeTtYf7Q07XVuXvI63FmHYW1Ljj4WaIHqv1TyPXh
PNQR5YRbeOAXHV6y4M8s+ckMwVa0dgCmZpSvBy+XUiyMR/PKkuI3gwhsna8twysGEJCoQkXwms44
k9sS6F3gTO3bfPNxXKmBaNodhlPh63rrfMufKETvHZEVfcu8zUjlmz+kGkb4gR9yfda/yZyvGCAH
CYQDgeO8rV3RdYj6aYc8K3bLPXw6dNDN1Zuk6vPW7RiJsfwT+IMMUE63AhGPMs/g+RZ4KQiMmuBu
NRKSdE6pI2Yt8elAHK+0ePdZHROT6k07heFIKISnrr4WFqLDNBNSXwmvQamEglyS5aBR6tNDL5lp
Y5Fn5YR2I4LS9C7Z1B789H+oh8+HkcjiISLpLrhcWqvhXL1kCjnAbc6BYVn22rM4eGKvAy/Vq+lf
4LbGL6SeWjpohqXUVY10DBBJWEiHaXZrvfnrZ6KY3IMC6cMXm6Fqjg7qmllDGFULKuVaLG8OE6RQ
+RRtx18BhcZjDCJ6gDXZfP5C44KDe5AEXvi+EcCBofMMHGJJ3gg/v1umoMgC3hJ4g1ZjIFgvhLPu
LWQAT/USeHGXY/kSaC9yj73BZBzIzmtZelyXEM5+DUw1/IK6R7QftOkAUtPOVY8gqswhsoJyUPYY
8AAMCmMD73ffa3YeVeLCSuSKHMI7a6wNliT//+Fbs8UoQDFmpUfW+QiZGKvaImhl+XRqgThUf8Vg
HGhhsZ2+YXHpW6bjrJ/nP5X/SlNdlC8VXK/RLmwwcva2y1j/0P/GYXj8dpFNBF+6QKpgnA5yqQEG
4qBZNOuboll3eOv8Ah57qCgnAf+TaF34Y1ujlJcomnyZcoUqak8tVrTzLFE/fMFIhA4mkkG0MY0O
okFDZW/nuwVDgxlWZK4f0A7KKB8pGvhyW124OVMrb5pLUvT37l/GfgwzyAhu3tLCJV1sOCTiaQXK
T4lwJjPElQ2ny8r8EUJxKh5d/BVcMiBUjLXOvKnKew5Jj06svoIAttL9KTPFDV4ZqLUDna6liZ1L
p5d6E9P6/xVWnN6PhKpNxBGPuGeMtH7qRwcrdggmcus2pkezBJFJmYrxE2oYHaOeeWdO4EKV0F5e
NFrfHWT2xwlIh4MKAGcbtklfrC3KNLFGq8eOUg+nP6gycFPi2XfSJw10s+gmY4/MPn3fJ6dVe50u
AFXe0pEJfTIJqe/K05uNk4JBeDgZJcE7B2e7YLuh2B/3TYgUh2Cn9cHJrc2jM0mG6AzR3EFBJhn3
4tvsFdDNlQVtCVrpL3zIu1VgNVV5r1Wp3BIuEZrnXixe32IeaxgU4pcIglIzMww5d8WpdtbqhqPP
Z47ieLpLN1o6/iExLVj9aMcfXI0upIFerhLv61WRk/raT0DW1XVatsigggQGbY/LE5yy04QqucWS
P5RtW16+CCosLKZbce5eGbMqhtBEsRlbLpXpJN17FQ0oyu9Mx5JLm5QyOV+eH6fM5vymBdjq+jHg
heWlGGjMo/Q299AvgI/JcO83TK/y8MtQkiwe35DXNkQ2aKBoXfTEZTTRTL1I6zoGp+0CZODfNbzp
MWCL6IDOTVIL2NasqTHC9OPVnW31/XuTqpdmDMIkDzbogJ5Qnubf6g6Z7PnrU1EtFFedGtD1XGWJ
xT+tdzNnp1GqP1ZQhedy4B7kj6Wm1JHBLpZT+W6Mf1E/ydgYy4GgsKYbqqeEGSzwwFbBpsHV3hY7
fWgoxwfMTqaVlVk1BhzX/kkkGuXKX/nuXa2tBrP2Wbe3Zjcu8AJGxEeCXr5lzN6NXHMAWEJsbNpo
5HYMYR5SdC/uF94fk+BdQYBPZUyXsD/InKFVJa662fh6TbHMqNHuGBVCYuyudFZEAMTED7lAOm0X
j7amWIl6Q/QDF3FwWlwc3OH2LwzSemYXF0TdCmiOsizim9HI+0tWBuoVGjMIC/O6O80s0nNx+srC
vA5ylY1+9YYEMa1OVeI5ou/DtFjqHDgiAuz5gR7zpuiceAsTrvP/rM97S8ElQ0+P1P0T8OFlpofY
fRh4OxTuC+sxnUeWv5byd+u7N2gJ61c/ZOU8wVDe+dhTrIiQw3q7V0gwWfg6nLRIlTxLOR8O3XUG
yp3KOk/HJ5OcesUG1WaUpi24MkD9dhBId4BDSUuN8NHw/6NTUQBNJ9Tr1RQwJv8KqcdjPlFNN/M0
P9MW7OBAnf5c3UPmBVOuNZUmbWJ9JJbznJa7RIAIMwrmLoXmN7ICTcN0H0BnTrytQYsfNOYHbI7L
PyVo82LBTloCqP4M3IxHy1t8YGPjJncePoBizfy/QWqmaKt+FV7VI9myCChdW1o0Uda53USVZNvh
2/Ncm95tAhyZnFU3GyxtWMP4wa8rcTO7+cJCQRt+RpT6Skqynmsz3fAJ/r47aBOwX/lFxY5oho/7
RgHDqfCQ6upsaG6G3c1bJL1TnvDRoBGarxd9eFEW/fejv9lTv2b+DVXIQqGjp1vProRThujk16Cl
OFBA9rLqxp4C7D7+Un7QsAed/60FsIFmQrovhwbVDNflEseE1X0ewCmf3e+J09doGn5ZOgEIL2C2
ARgK6JvEas/GvongkhuiFJJKZ8GecxwfOQGBac1pzzC7TT6YN9bK9LtjQ7L70SgXGmb0V6yWzV+0
Fr5am2HqSddOezpcsSJLUOhSvlyK/nLFCec9O/JNNF2mryn7nxTnwNhr0HTZk0kaDXA2416Vn+je
vcVeJQe5pm66KtbNnONvq7gdlmhkCUhLI2I8IU96MHOJ2UP2qN3VRTkKerpuGRd3m76znRdgPW0K
Yu5SHOV+DiecrzooNGgECIquBbOm8OVDW+IxACWc+e/i9g9I6ul4EBpECsGvblIAY1ykGdovF1UU
39j0N2aOPpuf8Tl1qUqzxMkh2DdSYdWkmmTGt8ar1pToHByh4eU4mbwyjbuZ5ZMzfveEFdGViwLu
oFTa8PLLi4r4iwmsXnLkPESM0cojGi1KoENbFoEn+B5Qlt72Venqv3/EY/WhvSqlEPLwObxIg3lE
v8ZBa83ZSoAspAk6HwJRsDFpAxd7IYI5OcuLbURvaWLKfq5vvMeZ4e5RMOJTsue+DHGIbwyoaccf
CCN9HXzvHQiqf51qpgugkr8tX/XuCCwFUiQdLWPrWZdILWvB/VL7KHUgMpw8gg1l+dF9NxwbujGw
bza5AFSaSoIY4AldTlFIaEDIMz85pHDjEW2DtcwsMOgwmEI+x6aPJlhD1IiGS5akjebmAnLgsrcr
8yoPftZ9LN0qJ6wnmGxHo/DMpP9iRZqg7HMNP3czdbCLjP3zSmT/UAbJUAh5HBqwubXtutqmpEV2
aUe7ki6JxG6OETiuc2U55yXrVTPMjkXyMm39s7SHTps+sKCa6aiQWvfehlu1000Fy4Fhx9RU2AYF
RloeThmpex8dyaMKbyjY476a16fxp7je4zaiJ77RtQwuCe4fGoZtPs7OzzGqt+yPDbwNwpGVwkjf
88w7ufjA8LTNrUU7TtZ9g5Q/yAKK05szNOgAAuzQOBHIUYUt4g0nTT8XlyYieCep4SrhRHrwnJYl
sVQ1+DkqRXW6J9BeVPU0T5hkWO0K4FTofPEVBifz6teABjnFXsgVyrcnYgxfyd8tusE+4kNDXj+g
BZYXPRMARPBCexdA7ydXaItj9PBvXPbvcDPks/YWyNS7VhkeeMpKuKhHMFnH2Pr3E08DSmEkuJvU
ebBwz4G1CRjikInjHYx6a80GR9K9B4uNqhXU9mJu+iUHC9JMLC2nW5bna0925hFI7SytyxdXwViM
w0l5VRFmd9xHqdip/IeBGspMuze6ASazlp/RMc2tB6Da/cKyEnU3R3DZaGvqKzghijaTAZbJI00f
/bikJjH3EUuw22b3LBOQd7I5nFz/CgPxGCTzLrloZDToHioIE1+OnIY12MnoLzrDngSSWsJHpTq/
/UJEE5hm/4J0v/fTqeHkciuCr/i2NOIWWutvL4rjCitt/DsiUWj//wnAfEotpuRQu1yNV2qzV5DO
/0OIWsF5jHcDJw0kMcLG3GbEQ71NjiKlFr0ev5fpEu8X+5Dv3kD8YlSzkD3cpXPc6E1is95mW9ZV
yxVEvyxb94iPww4yKhuxt4FXDd0sIP45XgwsTSf/K/4bnJlIxg+2HTGx8xTdTjoS5sgYV5FRJ49k
Xl613d9tBTmROM4AYSq8Z9ZnXYo0qGlKlqve+k1IQElzlDhDzNudQHvuBKG+9vk/pCuSzOuNS/2C
SZNA7RKPG7myOpuiPrQnMXNuo6PrkbE0HWQrQxyuSoWD9dUjL/QjW+q0sFHa3jIBYN0P4D9YPAPd
NpbPNBnxyYyTVLPngA8V95eei7nodxIU6C0xTeLtHWhsG1It+hNohdYCx+UqUEWeKsXJVMvFFVW0
qcMekBMBGyKXAA79yUDq83HJCtmrNjUg0zrqpKYxf8rp9bf7ge2I4YabwlDvUlTeuai+/pVt7fpk
LWve10Bqr+wNBBjRubIdmd+yMtNP6O06LToVglR5v1Ch6DLt6v+j9PQVYic9hxJ+bWfDV41h/htN
dHMAJBBisnUAJgCOUO6WNdnlDZGsTbq4otW+cgFVR45Fd1klmdSHnHa4k0MBRdFwOQb5IL2AOz5+
/Ro9dPPLbUn2taD4HQk/NapjPnh/vL0PkAs4ggdeHdziNXwLZgDFo6TN0ezKRI3oeyV6LaFGEhkY
RUVV1x8dgPlqtiC5mt0FXPrEGk7098aUc4awZ1e4DSap3/y8cjudivHKpF/r9XTsgirASWeuAXrJ
6WMLGwCdH1Kgmzwtj7tZNaS45jxmwJIb3VTqMkeslq3eR45pS+wZIvCyDvvN9fGuB0Z6n+05PuWw
JgGX1KzplBBzxOG5ahQxNv/QrBHwBQ3CcFyVpTRilArqJN3pdVl0AoA+d2TvjLv4GFfL68hAE33L
CKzIdeoUT0i1Pnr7drZiXjWCEzi5b0u3YldG+XqU1Q0QMOG8zQR9Ho+4T7KljFxMX3EYxMQ7CEn/
L/BjpYQ8VSA5xQ7YZ6HiJEZUT4TuP3BdpaLDWMwejSRyrW+SZf2k/8dom9hElkf/cigp0U5BWmq8
p9xdMo17WvvXevPByXSscyPzWbWqRfPR9Zz22jBuuOAk+AJT8RllofuFpebWfqHVBl8qokiCbZKp
UjPKNuckjBOUTJNnw4hOEtGedM8kaX8Y7zt766RR5WC+Ar97IEUDIfcm2o6bbd5RNkl+SUguBi2p
bptc1suIgM0XNFeh9qK4UL1Zp/si7dtW5f7KEfNydTdtbEK8IHubmPPgfk6M2tB9NjfSpDaBDrrV
PKxbgguJbWxH+8bmILiUdXTlpdhtWMqFJ6LwzAZZCWT6XGSblniKRjWkHpCn+uwNa7XFfD1qYjAA
NeHRcoClM3rKIJ2/0Xn+ejmqmXnKJq+wKR6ScaR9dGLzL/Fo+mW12/VJm3oR1mIE7MjHp40orfY0
U7PmCre2JSHaSL51Kmcf3d+vRj2RZOXterjgk42an0N5Zh4gcteneTMO5WTJsg3OtprabW4iIMjZ
l3f/UofksAzQWONuiohf/NGis7yoCYk6KnK+nGeh3pqaJ4H6spQO5gxgbpKVfFBlJywbJzj7G88S
sbX4PbacVxXWcAZpuFtJecvy3YDqFqr+Wk/RcL1zjMG/A+rpcd3U26GmLWsgmC1nM91ElT4zb7HH
yFl2tc8dybC8xirt2KieTpB0yAZO5tovyCVeZ4e+TQmGswg0yO15jNRksXpRuo0SHlEanHAjdG+J
yHjQHwFZxSEAkJ3Sk1TjJ4HrG2wpTT7Iou/TEo1Tc59G5oSbrvzTb0f6UVBs6b1gz3dIfSxP7HLl
ceYuLBNwuqWjTDsmFXHpUB+o2+1d+hWWOhfmFXRm6FcBv72BMOEE6I6NzcD5WOqiXIF5+51JrhS2
FSR3iF03WTwcxXUdnxBAjKX0p6hrOJxuRN5tcOqigl2H8Tynd8Gj8aLzo8cbpPpVFRvd5jcvrP0a
nIQlDVGqtRWmkScVC9i9XzvMzOxbr0W6Okdc2Apr+DMCb2ZqD0f6UOLEGdwq47UiRWSFSK2rCOee
RqfwnnxFsu4pc+hMU6EDA3sEIBnZUtwLsEBpzSQDaotnChp1uMR29TzaSAcT3GMbB8Jf/BGYtVgh
1mBSU4Hz3nj2Epl36Sanca8ODP6eHk9Oy6wk+YK5SZGXaJJp6i0m7NjBebPB2hLY+soGZM7DGsld
k7Lg8aH1WLMNgR5SiyH497TtuvZ0QgY/U+HChcPLZLXh6Cej4hpm8gsASqyS5/Fjz9046kvJb/mA
Mtlfo6fSpHpAYs0P77r1mS7CLk/8yi85k0jtTzY99/fZX6jDoVjnrPLzAU1w7Bx6KCO7NhN3anZ9
oPHTyMliOlWLBHrlsIFXJD7bC/qKRPREt+FvNf/GBHCy9MckI4FxJii+4dKHa7I/HMsySf3+gf8G
32cVtuysB8vY3WdDqCX1ZS+0oIqIulEsa0w6F6as5MCeblWcnUeU2QPiu0qtZi/koz3FyHJEjQrv
cPhwZgmwXfk2UtoxphDUOEJiRNZOo1m33FzVg2g2HQJ+RQ4zXY1ZkLEFFnFbCTIbakYmErY8dk+q
VOf3QbW+98Vyi4dHe53hfLIjbXKgHySFnFyn1hepNyNIq5qeYtK3JdkKNJXrXRelNzjbOzZro+NC
P7kGdHxZugy9rjR7CKuO8Ab27HpWzEgCJbCqn+hNqORahQK0zZixguiYWhG/mu5q11dsjjO8TVBq
G9RKkLKi3HovCjJu0wz9izXsUY0lSOinAZGFoua00TFCqpxLaSoqRFq5sRzWwMlnp/LAbIVStKyL
tDg56FpILG3ECazc/ko7zcIajsY+PUID+MyXMYyHr8m0/0cZmAeNlkyovHJZI84jNGKIfx4u0AHy
AYyzML25b3wfapVtI3B0saA+c0+H+SVAcjIJ9k8issob3tC3dAxWhOVRbsrUH7zQsewu6tM6w/78
7KSF8rVv+yF+QI+HiJ0qiYjKImqvvFznUyn2lZPMp0jJzHItD++Gk/qhyxlWwlCt7rcDHoJMsisS
yI5NOZ7AxrT+BciqjsxVDGIlROeHMziXh6apeuso1ZL02zI/SyfSMxcKhIWhiqmZtMV9pFuBFfyL
zKLz+KdXaypKRR1XigOVclu15Ptlc/MCEFH5f5kjXEAfOgpYFYaL4IEpiFtKQspQ0yl5WWEdnI1p
NK/ZwU34F1rhEOcGJK4h6W11hLhiDHFFCfhHU1q/hY/+vBNUy1ov0XtvupY43ww7t6LcTcjvP9Rg
7qzu+xgt84eOyOylSa1aE+pm00Wkvhx8yY9eVFcBq5AwdLnuDG6JwEuRvHboNWLnShz9j7RPXnfy
66KnXv5E9qYBO3EaCoPMNzjULHt5NIFx4XX9fr37R/5sfdsJtSM3x7M35gahCyamP1KjogmsX/u3
4nChY4i9Z82A4Dy3Nt1fEvuh3eLMZBZEQ+kfjmLZFJBd+Kg0jZGg6YW9IQABueLOhOcRg6ffOO9H
I92rlMOPsK5Czn5qRC6UyHIAOROc4SmNrsPdjr7rzFM0csW5PiwqFVQCovhsysOyeuvkM+dibi1T
LS00X/7ETmDl5IRYwCRRknP5DPgFdaB0eVT2apsHBg8l3WMzTzgxE5c4RtN4HCNSmdA29cA8/Cr9
iCpHF187qjdbRdA3Hh/hrJYh6P2QT6SrXw3Yv22GdUfNIu9u+OWGZihaeRvZeD4sIKbfPywCGbtr
f7U64w4IAujEj5UR6n1Bw3lcbdabl3o91l+Nh/ZCjsQtuf1Ax5sq06wJ2RqdwzIT9RZZeJmzO/AV
0lnNGGkEpJN0XI1wFsGnvC0+oMa4OTv7w5B+7jVCceVz55OBP6ebrTUL5X9kuHiH8cLpE/xQuEgT
duBBMBR5uicY/FN5VaPKB/KeSoKy80aL0xCb//KD3LzoCXBNYn4INKHAxrZdn8LyV1Goy9xpYRBn
Ho7D/eAAZAC1Y3WGCH7WY1IwAeRkabPde1Vt+F07Ph73tQq5sVSaGCZucmXV6KlkZM1PbUf8/bth
CcLoyTqX9siNxTSY5t7FZDcdyfgDMjiCKB7ubyeSRIHC6dBgtECbJtFVYD0ysYNb4Bf/RQNJT2Xu
TpFgsYNd8XBThmo38iwqAuvHiBx50U8L0T+PnNeV5DQyvWHyND514k5ArZmLqkrMq4biMBZHh+W4
VSuRONtXBs3fD61RmTeOnMzd5iH9dtzzeAghG5Rhz6Eun8Gqi4x8s6z2XUa/AGN72sCxhMlLvSJ1
hs5GpG3ncnhG+u1drwfXRekl1entKA3lR5fCrRQJbuyv4UXAcN4y5RWVbRlDya5ANslPltHGR7Hp
5OHDGON5HFG88byNgkkq6TQ6OQcWPQVMxMzJ/bALp305W2Rvohdo5CtB+HgSkcmAOC8iYOn03XvY
pM5eBRwWCC8c2fR9pLoCYxp5b9m77T68g4hP1+GJNtHBG560n5E4EGiHLbTZap3XGrZt/GKG6JGh
s5FNbkd5dC4rI3nM6SIfCvx8ItSZDv4vsVdBASuePXqIEKTplyujArBaR0/sh7yL9WbZ9do8Hknc
IAvCyDRwprCbI+Fmlr5SqyH0r0XFc0gNmB0VJHlw14vUEKq9QyoemnExSYxb5K1H0NIU3XklXXVZ
0h1tszNOJLmWmEy/9UFAknV0feCytrl1B+VIHZzUQDyLQ17u8gcIPUVW4qwUgo+ChD69eUpreEsT
YAPzzjPkCVbdctrTzV4BxAqRsonhzuC9b0NmWh777MiXoQULbOXspeAssiLY4x+qHd0ArUVKqnFK
mrk3UkTO9K/VOoEdl6oc4v3PMGRKoGIb1FayA/AmD+xHyHBZUGitoYH0AI19tUes5sEaRzx/1hmx
pvkrisIPQyfh+txJzs3MY5t2wUEWNVI/ragvczzK0cp68kbmKD9ayr5Yjqag9i2cck6yJ7LKjOdp
e65sMYP5yk4oG27d0Tl/TG6gDB9rkszOH9NN+1e2hxobEPlp3tnxP0B0EVJn80b8uRT9duyVNGAH
bIm0CpEqcZ7nQVLWl+jQRIVao9IBJ6LRFZcn9FgJaloCQK07u+H1r9htE2vxw0NZPcx6FJ205rzT
akbgNB64biAmz8C1tz1LMpm9szg+SCjCH8Yy+saldqvUk5xBG6juNbEaFO+pVWWVKz3HBnuMJCLY
PMZv6iROf8npTixp1W0IEpuofRY5TcB8BmHAyo/t2s+lU2dCHzlDNdk4s0SgRBKmcfs/g5Pb+lgu
flJDiyURMWSbgr/B5HlhzXcROMxeIAv+Ebcbtb3H3GISfi+P/rjQ/O6SqyIOo7nVIr3ohBTwrjzZ
4DVpZCZ07U5H91x+Sb4OnjWNYj0QJeqJ7UWYv52kfG55lbUJQWQNG31lKfAIWuRapYfGloRBJyKP
fT5EsSQun2BCDUjMMp6CjifdKTM3QvSuKB+7z0UyboqMYF7POl1Ej84WMqn5Mg/NT15f6XxawS2M
FHGbKsXtlcXzi2eWbS5qN+X5+vsOSB/3nxxeCpbaD7FsB860Nv5IlrXRYoVkC7lPYAX7XszbXt4h
M0Kz19WQ7cuNmif1dAYwHUn8Ah2OVTWD3dm1dL9x9H3S6mcEytpjKN+t0fgLIqjheJn3JN6vnxAw
s980GqV5wIUElYagZT1ORuPicYxXW/Zhiz/ZpHTEiAigLDG/ea+A7zqq5X/BWJqUzJ+hPy3LnQ2L
iu3VbD0DVvuXFJUcWxVi1Z3JaiG8gKc5C6tm/jFuU8v1YrWZasxlBnAWd2AH91TiNqbTUhZPZbnR
a234A9eql1vgKKQOztwhkAAaq63GliXK+4YN11LAT8jGES1o9UonjC4TAj4/LXNvz5b+5RQQUkno
AKMmPqKfLbWAeOJd3W7j4a038BLz3co8W5ZeiJlMB2VwO4k8LWSD56k8zIhrmxRLnB6BGYo4XTyu
KcIlbN551XEUMB7jTLnnvYw/0+xS1uzmub8DkmITAElt1NHqC++ZrLTHzHWPCqAecLHh+vSIkzPA
VBxn/4bcitUMZ6H79ufOpZgkr/maMrjwGFndjSqfWV91BPAfK3+OESspZ9NZ5RHMdXmuxNvG/pIL
XEgR0L1UrGIijParDwp6I2DrSeNXQlILiJuJap/IEabJ3JWbl9RwGjBXMJ2YCp8XIcUgU7LVytvx
4Hx9zwd69XfkC83VIHoKYbZuvgTLFaabcG/sHLJdv892Ju/6ZGuWCPTs8cbF6ckm8m4r7Q4TixkO
1gNcKxKaj/rPN4r6hv0G4cKkgBuUMVYeDELu7/F0EaTQnpmZFF8AM0dvwbOQ9NTbBOHe1pFaHL/E
KQViYqvtWxdJLMxsaAg5LIgQ6ZY00NmTrJYGUdZkxotdi0Xs3voLloPdsDlaQ98fnAsSfcHc0Jr1
82mGLDX5EYRopee6gLbMiTD0UvoES0EeNJPDq5G4EEWSQ7275chl6Rh/WyDFPlQ4gK0wwvinxsnB
sBSMWAFONsgN63tKmrAH6Cgays6hffrxhzLqd1CaTTXlv6vcHA9qlbjx/82rS+rtH1HYBdO26pb6
qxstckR/yRePE613kEBsRC0JbhK8qDiBUmxj535u9aQYfhwxutVjbp2gjTyUxLykME5IZTFM2ujw
JUIgRESpgjd94uqC+dS2PhiWvPL9WQ0izS6AZ5v8UHjcuh79h1pYCBhT5QqwSuTOH1FaSNwhTAM6
bzCZlSjcmhvcFnpBTRWY/O3xtFi2NKt67i28h8KwI/yPmm8mLGNAGGbi0TBuzl3udPdFvEMRP6wD
bKwLAK/dR0SDOzW47jlCz1Jl6abpeDQAUqws/FyEk38i22b+0lydUolPrEq3BjRaawpic14hquRu
P3Ds9jePgJLAA0FXFdGjN3jO/FAl3lNQwkdDue0vLbv2iS4xejapBYYZALgF/TMcZw/M2tEC0vpC
xTSrdfrXtf2IERmiLrVVn3LSRNK/gA7tLzcBa60H2af8+UDDlgoMutuKOdtScnuwf3tQzTs6urvb
NHIa99SJDbV6KSJsSm9iszmiPLFPTGZaM9abgNoANTVBGxFxyZGDKfRUDf1Vo+quHbJT1xHdi8Ct
GfUcqAAsTyALo/WLw05C0zPQgDmGNBoOaNCCyzVO0ZO+a6cIDsk/O4XHmsKPtHkt9CvbZQ7lU9an
EBGHK7rQP6KxPhKk0i+dAGqwd9R7R0d8fjHTuGE6D9xbUcF/JdQvnkBioSr3j196vn8RJuefaZa2
Mey/Ixy+Vv8PawXqr9n7ZRjuSyIhbzhZfEtSevQnBAGceJmySarQzCuu0ukMku/3tgKTIzOB5mm8
BhW/oYV2+txj4/DqSYmfA1ax4GeKcN2hFBo0xYG64bAQbf92gWHnJkao2gMiUJL/qRNjjRxFwSwz
GM3vp0qnLABmZahnyio1AniOk25wGrol3I5Dz1YtZdwGfY9zl3XaNUi/hM3mHlNe/VCLbuN9ah3o
lplb7a0RGXYbI0EmQk46VjF4vRjA1TdvL+lKFQWDk7BC/zPxu47eT3HE3gYfqFzX3oTJcO34YkON
M8KP3mOLGxNo6dkJdemuVgVTlqkYbVEWo+xAH1pCjoSI31onKFcb0yWlk9rjsMLNuvEqG3QHsBb5
Oizk3t+PVg7t04AGRYBekuvN7DDbQEMtZjbnKlb8zPtI7uoe8mXuIKl+xR8w4l5kwFp4Pp32ok2t
3BmnbgsdvWq+dqES9wuLBJC6bTKgwZINf8ajKtiEelJmDBlXlK05/qC9A2cY0vh/jkYURBGWpQ/z
NhflOwsV1inn4JLGuZmc2sgIGGarJ6S84ahMwqhmvY6TK7W+CtgOj4d4MsZtTkE/oRydI1MDlmeq
rDp52gA7zf3NHkcRPRluX7omI8SNGGViQ0FTXLf3cohZCexNp6o/QOuXmcIaysCC94S4X5lSmWDF
as5Pps1CKmmO5uVz1iocTwRsDRYEjmg00ZTBCFUgKTPPv6oyPjDWCmrDsVOmQi3OT7jqerO1XaZj
67cLQvHjUeaIyxDebkdGqH5pXKuIfRkhSdPAhWa2hflkApRl25FNDFf89REoN5cgUL7INcCOxzhy
tjA2P8FeEtQYKb+9S+jZ06ZMe7wCmTlZdAiAzoNGxP++RNqWJvQidVooTSuiOLEBtQvUhOAsvHl6
phFB38lmx2RNOCWAs4pW8a9R2YoELPwbHW+o4733ICINf7HAJ2DCWGRhxj6eRXJ1kXLFattELr4I
qfuBnoOSMiuHHQ//xmYoJucv/D8D7C3A4R/bBfNBiMVjAjfY2jeaPeg5YBrr/pf4HGkzrKRfU3fa
Op+DQwh5iztY24AXlFDSbYty9zkaoA9tsPjQ195mwhhKG4Y2UwZdWKnBPFDgZ2wjfyd/xSk48P3T
w7uVZqCZi12gzoe/v7J+hf9+u+C0M98sBSiotAVLDHQF4SXAcOmlndAxAcKxmf6Sri9fIrH0p6gh
nuqdX/sTBiYHjsHzZzstwiw+I3ryT09cXpaF6IhvuriWNCY94WMJhRKR0TI1puJWVv7WceEmhxe/
bSrE3ZjsZD8GpItthQE033lkQ1hRZVjdk3i3p9uiUvMN2Dt6sgytLKvZYZRU4o1rHqc30A9d3arS
LQGq70pDwmE/jh4EoIpB3zaVx0GlUSkBMtDgVvg7/zTFc9gLLIoj18SHp7sofj8E116PqrlMdb+0
E6m+sZXtYompkxt9QIlh6aNlaXIY3X8VpFEZFz4ePo9Pu+9LKVND98/glyHqQ5vdLSS5XnEzhr4d
AUUzo3un9Cdd3zdqLfHX20LwTm3JJmc2BQkAK7lAOjYFGVndo5xZWF9klr7qEs6V512tgGpsGkg8
xjabW77lmRTiohc0AGPLPGcrNETbYbUAaxPrgD/i3eKo7gdAnFL1aWYfMWLZvheQbAZjxKuAkfYw
5n9YL2kj4VzzMAeyMAP5SEh/CO0DH7NOB4E9JFoTu0PYoWUaBeNmA+ffC/34gH49qz35Gojk1ShN
83XD/pV18dKU21oU51+OOBPz+/9oOUhlbfWXcviLJEBuiQ3qat1LPtsvg/iLsPQrqCj7y7Oj+QKy
2Y08ni/pyqNl1R94WW+7bHnXDutJwQFdJGe6xAWJBV7mOwLNQSSIME6OdzwFeiolPX09OeEJsQlc
2n6i084BSMaWqICoieDZ6NRFW68fqAnp31xs3Yi8Bwok6vO4B9OzpMFBdExMroCXeAaM+6q6jJXz
CbBUwIM4qsZjou5Y7rMxX+PApJ01Sw1yTZ+5nVS6uwM1eRikxkruYpZM8AJtf3BxNiOHXkwZYbiZ
y2wSz3HPF9ZZQBC4YIa1TCGHUUnvqaTX5+tsI6aeQd1DAAohA3G/54GHIdqGuIORQ/ChzWduIF2U
IMiFrKproUMeyg7lwV2J7tvDIVwv2kwk9vhpqFh/6kaH5JP5j+3uc899gbCLFiaExeRkZ8HDM7Hw
f4tpH9ehm1FOuobFY4UxcEa361rYTM/xUT+cS9XdGLU7WXoNDkRvFvP/RhJXpjV0QolFh0gr+8bf
y51Fnx6mqSZQP2jV+KC0UsRtDzN/bu+2zXnuiWa+nNtrVYT92Sc+5i0+hwk7dZ2iud2mlOvFbJAG
HTzsdrY0q3RTkeBuEm4mL2AuwSl6Mbd35WhYHOBcokuUIx/OnO0KSgW4YeV69uD+0xwv1ticM8uq
Lt3xpbLm5uWDEa1nOFtBd49vI8VCxVzyYEBfkoTSxMCnbvsPvy1eeNqJqNB3Z+o6WHncTZfa+BQV
/Bq/TcPTEAWKefVssCTPVocbuYAE7+y3OnT1QEJx6vOBf7gaTexmrg2q0UaD8fsbABwh4L5aYvfv
sihouVJakhBAJHu9tzICSTRgphFRPMi+tQ47YNacJBVb74F3lf8ynlHPNVC58sL/IEzzNdExFRiO
qf0nqRpFZQkJK9QG54pveEJoaa3+SO4jyBtGYqdvnz1743qVYdq7cDs98+i8rV7Wq6T7o5aEERd2
tOaC6AqSx7PoiNEvcMLSvlZo4ovNinlG4DX2sY+4XaNfDZ77FH5Xr9Li9BhoS/XW6klF1atFCrrc
nC0Px4eu9M+WMoudcAd+ajPMN417cqBApOhntkB7670myw3MHsTBt8D0Q9VnuHktCZS3nZ/8fY7X
MSyVwVwOesqG7PR7dbKZa8CYiw0TbshOerLrn7MZhPLxMicjGZzNrgqMC1fhGu/1cxm995bKFfvK
ERx3fC0pyq44kJ7fLNZ1HqLkE0Orep8TGA8dOwLFiZF/7hQ815yJsNHnpvvQ9KbBYrBpgnM1flAB
/732XGelTGCatRjAxTxK8v0B+2NrDDNhqvyZeEH9njg2GxibeOKwO5i+kyYPOKDFEjnU88FrC2md
LZmGa3fez3nJmuP9/i6fvjpCNTOguLYgalPl1KzQFdKV7D/q2I69bHyZo1GemSVr+jivBK2msKh1
HW47Mmwi+UxMXyU+46748Qy9lFghnqBScF5HRixHC29xiwFIDJNQOgkGa+A8hdF3rQe7pHU5EBD6
OmMEo91J4OxynLpqamQ1AUN29dOp1YHNuX6tHt3T1F8rGNELIRcE9a0u62k91mQTWcePE3sdry2M
LhbcVugzoB7g/vPxu4GnUKwsy5GDuqfPjTd3TQmAk/oDPR9JUGYvhzQmhb/mNES28WB/w7IMYL3b
SeDEFCvFPgPKrNxmiaZfhIDejseMCsW+/LY7bJ72vXflzHk2BOOY7jnzXoqU4hOh1WwsXdiZAZ4J
A2MATxSilvmpTrV0MCVleHuemHeoaDryMKuf/sheZ7Du7zLPBLjh0Y8SA8PZ2JynjWlPwL1dn+0Q
C4GVkuB+EHq9vuCWhxmb6RPHL4bpvAtlu3jbDSvq1yYa4phqDDEU16b5TXRVkgP2SOf6/8RjS9NE
SxLHmEDPlSVXIUOkXeODU4mDRjVWuzyCeQbvpvzunX274OMUYJDZ9qwpeBWL03lET5IA3Iql4nUJ
uQexdHo60cTy/Ehsn38YSkoroCrQKngbyg5i8TIvKTZvc83hhEB6W6YK92Z+WCzrialLreHwLbIq
eud7alX67lb1Qlpn4tU7WPY/0aNOrOKxEKONbA3rmMRUD25CjLNjOsT1vLDv5F5OyMY3aqgcUs/u
mPMhT8bC53hC+WFlwW2v7aPrI3ZgZU8zVRrv0M+t8aWCfO8VW+vEkL+ajCVJlgOwxsjhHsl7/Rhg
J15uBiKb3STpiuOJchSNGA8NHWJG2ShqgZ3c75h9Oe39csaLmUgX029fM3ug74pLPIsk+BMVYg6W
FpCUenmRLaJzpSbPhBwFrX8SgH2PdnBW7LoHW9cyjgyS9/BVf39jBRezoEOOhKmOaiQLDliPzHR2
pEgm6/kn2Q9gs48q0Zj8X6U8l3fICFvogJ9rSYPDtNWSPaua9VEMuui5U8HinXetFGt+tGljC7B3
Nw9Lc395zrrPI18hxVbFOrdiAz0d6K+fdzHwYajrQ+Wdupb4jOM99y4VgOQPqEBa3JD/pK217bym
U6Xna5JB6B5Ov+W4AZObSTn9mRQNtWDxnpaDMQTbSI9d14UtDEj+qubuovsGtuQhtavAjNsBz5DU
I31EPUrmKmTJq87ro2r2bYYkZo5W1OgvrBtxqigMy3t3LiwKg7p6NAnyj0MNFcOho0vIOWPj/Iqr
2f9JF8A/GAs1oDpUP/8ZV8J2wDdpVJDWGTctk/rRASR4QL6upJMnG4sweT6HT+qeFr8v5gm/efWL
9fY2665QTXzkeHCLnd0fHxcGFjajzJ5NrKxXEwrICbKLVIjFCiEalhCt426zGX8o6D7ddyKQqHFr
VKZuOMs7g80ZEniy5kch88Xc5i4kCdG6WbGhB5N8nthqXv/TmHG6TIbUkA9ki2U2iviUBgA0LrLU
oDYyaTIl1wBZsZ4RwSyxvNEWdoz6DmCrn+IqWOfNR4J1HWC0B+ELbc8VbStOH+sDRPISZ/mJ+v7W
hw2h76vo99XY91HmG7lxcDgf1RJki/XOkrdUfTsV4P8x/pfIMU4JsSVnrHId5LIixpy9BQ3Et9oQ
C9va88HogDbselLAu3bGTG0C6E5yhgXE/VjU2Oj0aA+1Ko7xoOuG7wIjYnKI6rkMjWlGxJA7z19B
+kgIMs27hAtyOuHyujJaGUop3mCu2tuHO6ztmK5EdVzOc3jWTC1PuPm6N15JlEhXDBRCJVjB62Hb
qOkIdY8SZM+8jbeKvyuhqcIuGTvdU2J8oMGa1a/oG80WhkYSAASpvHDu4jjIfN9PAJpfpXBpGbk9
OYBttoBSKD+54gbv6fhPa8ULTk15M8DvX/s/BaG4v3l484CcGZ94Tskb68FV5a+43IE3U1Y+tVDO
LIEG6wAtqcaEwevGfECb8MGzkl5XzY/+Rg0DyGgUZAu7dDTdYDucpZAPACOIzaNXw1F4ghnluypj
7GEiuDgZGkdqQCIwrb4e3s1fdM/FGnaYKbZ3SO0vlyMTyVNTMJN7lBP0aWZs+Nq4Y+YyLtQoOiMa
Ptw8/rJss1plyajp83Yzx5GgFnRML0t6LUco3yqZWHlv4B0ac5lq1MeXmnAouYcnd09kZIptk7Ep
zisLxnkFzpYuXj/+7j6BSAQJeMV5zx0DjfXn0s+kYE7i21hME41QN/Xa94OddU2ae910PAzaeG/D
PwbetCNIK/8WEFUXTy31/lNI0EV95QYKx/cV6EJmGb4t7XobjmNkOlIw+d8VYyU6YMX2bHncMlAD
ORMkTuh/++P0RGLYVmAkZjf39YS2hUVFq1QU1M++Xtq/pCY8A4vIxsvLLNO6KmrzzENsNFbs6sPR
/ZF/UNx8G/zttwJRVA1l4+d5Wo5flO6rHBhzjVAMksLatJXTmkGQrc/lLiBDsvBpZ8/eKLRIoyC6
NJ3KNoMnPOyLijf2yP+QrAL0ZCp+jJFGuAx3JjBVpbDML5H43epO9I/ZNaxvwm7X60JNC8QFs+Zb
+Rlvhjg5ETuXtEWlGOKlWsfnQgxYQlOxgsibag11OkAGfE90EEBECTxZsqO+4rtR7z3s2zxbtneu
ZSSx0B/H4qhDWi7UEElvw5LxEnlU1WeIToubP594ZJH1ueohpQkU5Hi18fwipyyZ4uYN5oyZmDjt
nJ/e6dI7kUHIuk0qC0voBC2S+VCR4JUYnlSxFDiXT0ksSIO9hMGGrHh351aJtAsJ/gLNO5dvqkJJ
r0gZiiuHQFBcP25Nb3MH4JmpEZ8NPINNhYjRkeMbrjS7F/ah5KYQUH73Bz5cRlxXOvEZlE5Z0/gz
xOJNMvIRmv9jZ0/TKIiaOGS+KnKNmzzXzY1xoaN3qYD8lVn1Mp9ezLQZ5vJ4k+HfDeVghralyAtJ
qnq/Lz9tLDgwLdjtfqR7pLJP1KQ2+HSqNaQY/oC0MNvqcE2+L989IzD5uD5imCEF+LdnboW6oDu9
lTVbnRAjlAA41YBpIU7ZYeSi9p6TIM759nUIBq+AJ84Ma2Aa/icH6DxcieC8pyI6Igs/z7e/ruTF
UZESRy5+tLJPWmeIZdvpeKg3PjOxclFPynLl7/XvO147Ual9EID7fgqayWWxiktWvP0HmM/b67Vw
pBjatNww10ByiWnLR24JP40c9JIzzr7t5aW/s5cfXbHwR2GrSyugBa+U2hb+g1v39GOaQvkzODtR
oivL1FYH44u8KowyupJW2D1WRccaDuKf0gjQlpMPAVZyoGILvWLPttNGEUja7niTcDRqJKX3Q4Tb
KB1xIYOKJCRmP7ORKuUwLJxqumEWyfFNfHYZ4bZG8pAT9ejHmrXwIbTbmg5PslBm2do7L59v1evj
0pT4aRwJdaVN+wU87vTTgaemtDwqEQqx7qTWJJCWWGHe+GyHJtXZO2THxe+gimxGYmIAUPnSp6PV
DuBO/v+tgiY7tHlnb9vt2C1u4wHwO5GqjtAR0rIijC04TDxD9zRgUkWiqw2CXUaR09r06GN99ETZ
JESRwgCS/+W3vx799ijSKLjpLsw02ayQxMwR+fr2Oz8Ih8W48NMacuz6VAcSPb8j4Z+e/msZcp9U
1DLZq0fyJ5lBdCQnV0eW1IASttK7HhxbPSCt5hRkRAxNpXD457ct4J/f8z4U9DdgwSTIh3gd7UE7
aKGVEFTYzkCgd7l4AINYaQ53t+JfvDdyWmmFVoUeRSaLrkjCPg5zunGaJ3cQ6y4tlBFrYP66g5Iz
gNxTe7DxVDwVYaaxJF8dBjyRkBrGGFf3LD4jPbjZ0afhmnAX7rMe9zTZzYCQuUAgkMXX3f7nHY5R
U3wFGdmx/cHw5U5TatuVpeYFWKKmxv5NbTUZRKjOVg2G6QqlAjwqdywEafIVe+f4ne3gd3cz0igG
jyVMWHCqHgSszi3VGmn5AaHe9p1sIseSuQc287PMLG/CK8SGR3zG1MK4BIiZrz8Z5EHGYdbq3/Mm
l/2DSkKIsw7C1gW/Zfpz1RlzYSIeGSvOdD7a49CR/jKIoookZJlrSqFmma5LkWuiaE4CnJkUPfmM
NRZEDqMdVTrTey+TJEX97zO0G8I9tVD12k/zKQ4omLzF2rXmX+7sQdyEpzfTWpOqgD7fGikP2jWB
DMAd2YgrTyuHurD+YvFsWw/sd+szWw0vMTlllOX2YtpVdhgfKXZ2jC7oiWHR3M3yjL+jl7yWLbtA
LRy8MMvBLYejm3r63p8X5IuGIBROic7MfI7XgkBdQAZqG6QDmg8fn4A3uvjlhtSluhvJHTskGKe4
slhVT1usF5QHBYes25XHOGC3oKwauZNL3GLut3+UVC9oRqMEl3g3BFGItse3LW4gZtwf6kfWtdQ5
zXDti/0SfxcN+oL3HsmeQZXbDaswoCc3rwc8ycO7Y8t2cqNAj4J7snYn+jcuONTHTQ8D0WWgF3/5
jq62nspkPfs1POuQIhIqUbiXpiJwXL/Bx750JcqSAgyZv8id8fSIRBEq55k3EIkMyBoesFBwVsjh
VFBcnZXxcIPjRTiorPpSvjYFqj99Z4QhxXlW0mzIRtTkbQ4sTizbuM9nnxObKX6kCzchC4FAp0zW
uqgxiNKgGH0WD5a97Ctt+4BOnVZ9j64Wm/yoxPzX0jkA1F/86u7FuTFswWGiMHXw071Y8W+DFMTu
gspnySZtaQxWu4EFX179ErMiv2LKhCERKtyt09KJ/3pI/s1x2UB9cn7c9RqJyfHxZ/XbVD/NHmG4
jvAcBVXtzI9GRqC+A0+QA1tBaighOxbaLQO2wteHXuO2j/v+5E8qu6pNb+5ONV2tHa6wXVTIKa/g
EWU/oF2GUZ/moNkk/wDwLRlPxo+r9upyyX/8eWGaYJcY0uFn4wuKyohgsm55VEoPkyVAeBf4WVjj
tdDUkmCItOmQMS+fYTV7FiSL/vF6EyQTyE+6HcO0J5PsEcqLwaDkd5MKGv2VWgNNYONlrl9X2Upg
nJmMyTGkgDpk8eXVFb/7+U6JzcmfcxBU5aFS4lh01DYgzS//1If2rlLPkYabaB3HwLqwKW1hilly
Oj+5B4xDU1Kvs4tFl+3YDyioxqciYz9xUiHBCWpsxHcAiXyGZ2t6Eak11ZqlnUJcB7tqUmQy518L
VJMk3s0jyaMk2DBxUvwselc9mgFPP9ZKE7zXrg5QrU7sWIJC+cHVy2b4kJIgSW/cYedWLPAKOWAG
KGPUzy6nBu4ujbDoibzHkpc1oxSTlrJCszLC723tCl8ZG33J0EidQIko5r5BUD45FdKSHQeGeZ+1
9mbh4THVzOiGJUElZJNsFivzTgkZsoYJzhnCMU6sMD0xIaxowCTIMf/EaEj/FqG5XV4V1aj9gCq+
WmxP0EtxPjfyc0rhcvGFb9V4oFvnbaGvpPxIfO8+j1UmAC/SKv+gutqgSFqsj9PnjJbXHqwfwUZR
RbjJJlxY+IUlBvYVXhpmXs1qMOu8+nwMmfLnsSJ1FoC6/kOkyo7S8zEp+U+QMA0de/ZsNR6ZbLqD
HbnH2k60QNeMxXX5o35XGlEpYf0FypEZeajkOrEcXWI/HOybhVMYxtlJw3Vodx+Tyg0IWGkW3aFx
WsKxjp+5K3//7oUsk+LTYoUgN3L3Pd3lb11yNHSWGYuBhZmrGlZluDPZ6HDMuSJdVIy9KGSMpO49
m07IpGTtZszF4BShcsks/lGs0oUYBT6YFKj4t/Vq6VtcLcpOhpSV61BFpJr2CZh9n5b/s1HNsiv0
0sHWkB4pQTVJsG8xYWJ2zI2iYUNK+QsAG4v3cFFh8c7tOxlwxcLrSTfYBYVpvvPQnF7djsCXFo7u
DHDFyw26ZRqigDBYL1jZ5RlCmKtPQ1A9nnJqA7RY4ligWD+pXNeSMRSdfe6ZBDZwsVf3tcVoZmX7
e3dz4FnKnwXBpGmV/3aoNWZ0us5yxN214PhppWGAP8zRqdpQv6uBunGr0Oa4bSbiC4/P048o58uu
UQ1QXwtpMMlOWTvxvMyQW+UTeajsozfA4ALLnq9+OTgyvt+xB4FAmcLSj6g6QfL5KeH7yv2actzx
Ytwa49XUt+cI+xwXnGSnqfxx2blxak4GNNbfoE0YkKgah8eO3sLPnORqMyp9J7Tpwn9CyVlTtJog
+IK0f/qifiKUSFvY00bfnEYdM4xw7GtZb5B7wRlczids1B4Y6BmzPxDF3BO24FKG1XOJRkAJnKFw
Vzcx8Q8YW4gUt1t/uQ0xuZKQN0xdttBqs1pv8+haN7xQ2IYS0THeD4PoKhjazdSeccDF4uKAMBvi
IKMwtjkrZYk4539RlYiT/dug8s8zHGcLBdLVLbaBIXZOiw/850y62VrGKT3+qRoGdsHO3mwLWyII
0G+V+KnaySi9QgRUNv/aMp9R2n73RvYhwnHJhh0Ii1GEViV9u+x2O/OIzALVJaObZ/8mbdma59fv
JflyzsQrJJWR7a4iwlxr/rtPAFx6Mj8wDGjplOLo0UM7omE67pgEGg7sbSGhfW08EkysjNmheF5T
C4NsXsS3PP89SOZKICvDSeiS3G2jsNvhjidTtNZ02cyOGRVkmFXNUGa6JT9MrJjcByKtDYC3jHuq
k6l9XYZ9ri3faXv2PXXXrKknbysOoOS723vVnyiobTg98e1Fcm5qjM8AJICd8sMw2vjXOkiccv2k
l+CbejnA/GX5tT+lK2UfwIVpj0Q3yAJqHXT6ubwQWjxc1dV4uj3Ta1Fs7JCHxyTLGjVfg89duDhp
pbr1upsXlnhGVcWF8p2u8dXUaLKJEnVlnqk7U4hLD2uEBO2n4XvJBtHMXvK8aFwdwD6jIWB8StxC
jXxOVI5t+9Q+AgdUUaw/DjqyQwPwPrm/UK7T8AF2Woz80zH2jANOm0b/j1rkot3SdSnR2E/qnPp+
3EStFQBHSRINUrONtHYiSX8CQSca29OfzGFoHIpsQm/RelBmYtj1XhWDAXvLTS78VsukoS44kkxW
yiKabMvP+d0EqxqXJBnmHyEc0rhrnJUOGbPecSv5+qldO/JV9LxuUYBBwlJzur9bjHQiyjDC/C5c
A1VxisfApmyTwunHcprHDgK408R1uVTy9Hr8+s/rlhjHv/BOQDVzkxumY1v73NYCEXIRy8m9Ahy0
5KngArl7hEzGgm2+P5H2KCHVwdlStUEl5255V7PQFH9FzKt9WDTfoghMFozerJxsiEe5GCXj+RrJ
lX7O6YUugPp1Tx6ODU/YZxxCW/2ol8Of+bYnJw/CSTh50cS7KxiTrlIiQgJgaYWZK60UE5YQ0uC5
5MSZVZnseic33yQg6o8PwfHf6A2f2WuLD5IDxa1lh22dqgpsnA+OrlGjjbrQBul03kKk17161L4a
2OgyEwTIF9EuGNiOFJ6AVd1T+5jHg6URiwDdHL3+Vzs/71VHgc6O7lJJpNsU7A/jav3oYYhdG5QO
yPVB3PhviUqyWyB6PnaKAdYrE03f5ZsWTmOgwSBBBy2USTCUnMZCGq7o6+AVi3iyfYYN2ZLhAnCP
mjEDhY9ESSF7D42clkRJTH+2dHyRzvZTIhEV+eDIvxssO9axglvPqN/qy5sjNYBYeXapbcxF0Opj
eKE+eiLIqQoKwFI7ofgVq4afTjbIX1+UZDNXOuWVOLj6tMBrPcmNBKwdHoCTsK/mJfaKQt56oDUl
rLyTDY4x6ryw8lEjC/gfizRQkOLxXzdADp3iFg1EYuVwu9v1k0Tvsd1t21UZP5wKJEjmd4hBaY/w
5eOy6kzX8Los7cLlRzNpcOveD4ViGvrZBS28m82lqIiGJbqc/GGJ/4BMVUdIJnATdlsC72im8Nmn
EUeSA2pzLtqZrDprmudauApsdroneSTtbxzkrbXAJ8ZsE/hrawaHkLMShdao3SsEoSB2e2GdP4tq
BI9FNngS7NgNtmKdeDJ3MkT/yKIQ6eJPrATlJH+v055FJ1dNEcrp4q5whFq5dfff2LztJzgEh2dv
BwQwu+Nl2o3AG4yVJzyVUgIjkNf9En6E2KJ1meGzQ1UckoRsnB58o+o8t/wFOqvvI+5A8bfgIVCU
emo6OOVPw+lJMircuS+UcMPYY0pQUPWa3lu1hL7VxcaF4xPOHYcxIDlsfx6gm2q6s7Gag2sE2OXl
K4utqFyT8j+i4fLCmQ/8cKXNjG6DPfewdLhuASlzpueD9bevfNS/LRfTZaLOiOWHgOXLtwAd6PMm
0hbqBc1mPi1y3YT4e/XLLtTrGAffNSqZQD3onmsdehEK74yrrY/t1Nn1s+GRAwGUv3kTVE2vc0/z
6VzmlGT9+tepoowO553cESWIohfjCaK5Z6O4fXIdVaQ2yz0tlXgD0UfYmYcK5cvRdRHPP6nuGLLI
0UhVh8tjYsN2HZyFD+3Y58uw8GcUTCsQ0fDBWuiL2ctV1M9APv5cC74ZhrxWrCNxVCghPUXUVq29
H13qlCiJQokSokb499v2u+gU2MeD/USOE1wP2hN7dZCaIv2xfL8ZZ8FUMZKOGkOnZqTW5e3HwArM
3uDefk7zEyIARw5w84S+BVUG2A04Mko2jooscatQfq5dJkkvHoFOQcHfIuHI4xmiqAUCVGeXQQPp
cQqpPGpRuqg1hRUVCNxAJjAKK5aP882bhouaxKNWz5J6oYwSHGML4gWST8GhJjunodk1hJ6bZV1g
T+KuGwkCUbkIiKXHdIOhn6jZSWJ6Bi8gYWrkaIu6Rd6rF3ny+zx5srjA/C1vXtA3OkmOVj213PJJ
bdMqAhCo38mylLqRNZv5GeOxIhDgWo6uIFYIwd0DsZvLatZsxBV4lU2fUsepEP4JiEgU0l993XF/
Ra2m9SjsLyfyfy0diZniyt4WPFevKlEx3DSctiHVMvlRPDW6/LZbehmW5m3MXzzBO9XH1cAIZ2ZI
XN7UHEUsqGnvCvhL1H2/umuxESVqDGiNvzkPgwFjotfsUa5AuobcbsypSewGPprRwYrgofv144EE
csP8US8iVU3CfRVmBbcCoObTxiq+bJjWj1/gg0TQvE0AXPfyy4vDx4195z4ZlHGH/L034oGW6yzD
BXT7L0S08aRwAVLBr46gYC4W5QKwyJ4LAqm565DXResCSHd6gqDQWaM5aeGN4raq0E1460SvH2zb
qzquB1U/ONJglblB3kcxyq1DK4tzA6sPSYof7t2Rfn0zIsRyuZY87YFNtAAI528WTcSqPX7FMcXQ
1reieLQ+4xdbj51DGf7fvz0MfOpC49DikqR5vQHfUj+mOGhqBKZVPBeaxLitLKOOOfAY00GhDtfM
QEcUebIW43UplF+QQzb7qGfx/AYzvI6R6oSfOMouhktSRML+GGqEU5+lxNeQLWlEoVc2NXRgjNP3
qG5nyc4dMIhryTUJNfC9k/6o715Feglfgc3fKrAhoKPM8V0mqrhqdZ6bYKRdwPFNrhZXOWhTw7WN
SJM+KMs4A51YrZTlAwOsEI9vWDbK7SN1fGWuU0cdThXIpJBiYTsG5tCGBa1z8zODP3nhSciMPkEw
Sn5Hib16QK05MRf+V0R86ONjg4MwQiNUonMfwU6gepARBtXJFJn0Br4C0QHn4R2DQJJEd3afSYrC
ipQogJJDwfPs358Vxnrg0cTKDRcKoWksYaqSnpJWSxQ5lZx01si+hbM6073jQrthYejA+2S6nI2g
5iBCRNPINM/dSLZrMJtNPmY0qEi+fV50NQrXIF/sChpNdOkdMOr5yvUgcaXZdgmirS/Hdo+U7I0V
WqNFHV2PBwL/qZVz/ikg2hHnoHWIjfy7YhcEZ2pC41vFBO9NeFG4BLTZoMwSYtICrRAlfo+Ldvur
WMaxomrsJfjhNgqvONU2tU6Gal9ZSfyqw5K0tD0ZAJ1I48L6axnwYs7jbUbwo3T75bmxQKxxwzGH
f3MvKP/BV5w472lJZ84hguamMVU0lcwNi/ggjyqwIbHE6wpDUsOdDsjz9qdxd/lZjmTaLjJtvvE6
pFdSFjOO6HstR3RznyXO31FxPGZuj95Jgq72KcJzzpia3uWPAH/9YhjP2DKqfsMUoeJFPqP2+oNa
5e5TPIYbJ15oT34iLFufE8EJUxE7VORnPiVP1xC0cj0pUC12da7CPdsGIyi0IzCABSKahjkdiABm
wlifDnjN009P2wQ5XPfXOSdFsX01FX2Gl4UKhRsv8VnhsPaMJ7KPGfNwf1QWKMM5z21lrFGbnzpW
+RRhpMbB0OCQ8rmCACLS1j4yAtAtDf7iMk4NPyu5nVj5Js9V+b82Ovf827K5dnh4+gMMIX/uthM1
YVszJH9TdUvL0sZ26s4mDfc9eL/C0vF91dgb0oCXslwWYRYiX8vgrtibXymvd/TNzPByZ2rYun+y
rOt2HFVMkWgZgNY64ztZEXL6RJeIGhrqqdF0BVAshv6SF9xcRq5jZZSCOFPVrkrIw1nm9tjQDpjE
o/9SmKFMQggoHSCl/Q7/M4dBfz7bTSe5kH0UngmeKdaeaM/u9qDAN+c5CzWBM8x/nQRqbgD0n6me
+Vbju0yfs8qvasvC4eB1R7YpnmTym4+TXbVV1j6pJDsUgM/donqgdz1EajDnXXSw+M4SAj2IJgVT
UaO+UgGjTQbuoBw1BSWOvWbV5vEpZmxVyjjFKr785/Hp3tlPR7Hu5dU1rLmZlTP11Zy4hxMkB0ob
FFknSzxm/RFZkQkLgOsNHjqFTjgtzuZqeUVw4cdcISbIZbq36RXw+tpaq4qHB7ovF4OAb5FOtsJf
v5EGC8LrALFkbnLAxPIsvwTwvuoUsZkrUcbWkQ8XglJ1gfHpncxOaqa9bM8pCb5XhjO0nz5VLXzc
UdXcRMUlCsOgjhwqJkcUj73gS/tCRQMTN7OD8SYBpO52J6oe5OJue74GVIlUwpfFq73fYGU6MDsq
5dUuvCTPfE4zqEsbPqxsWb1FRJORTOz9hXav4l4utXbqqVKzUXSy6mUKXYAqDpPF9WWVx0qnXp4p
B3gHMC0S1A+yW9yZLBGdB4J9VJNTxo7NcfmrRthzy6xRJ6cveADrrrcbV4w4ly9d+JUpKjMan3ab
n4WJZzd/TSGYaPTGg2HWZazzyAASX5R4VD+FbPPFoWgNRu/GzIYrHNoxS6xmZVVlUC61S6539QjN
MhHbwLzd1G17xvMOuR+udmIOAKlZPmphz/fJejSuk1X/5ieQ11lSJRR3O8CBpbv1kkFElrLcHdJK
LVVObG2wwSTQCk47wgKhNimqM9hN8OI6FNiY7oaZRb5cMr+BoSLeM9n6740xhAbs0WRwA74koUHD
nl07HdR9G5yAo35KU+IeVN0yovnh+4twT/sSdsQ+tREIozPIP3jszd95UcpGEv7lv2sS5yVGGijy
YnXb1R38eVAMNymHSEuKZZpViow8Ulsad1ZjGDX4q8XYfW2K+cKgqnzHuwtkS9M5e4b0nRux3oR6
S2BqcYO9+MW1IPGJEB9u05vGJU9lM1/JH5/kyP+AKCZJc9xHdN26dVP6rI8frkYUh0yLNGyA6gnl
Zk74kWOIdU2Hh2zXmXD9ik6mVsVZd1Bc/R2QG39OCQwnRXdyh8M8J3S83+cZTZ/q3zanD09KgzVn
lKFrrYK7GidoKQ5EZjglnjga+v8wFlxRk34aogM2TxIhIqhnpPxE5V236kRP6+XGbGE/7OM56SK4
Wn7dKUxLzG12T/x9kb/u0Jl20E0lrVPJ98Me1aaWcYnFVoZHWBAUUzMvoe10r5tcnFQz3MMDoX95
jjSZvdhU2L7cEhIbApek+EKkkDcm9yY22RBqOcNgDiYWqo+Aj2vxFseJmsqydQ8XTevjRN9ALB+R
HJUg/s6/t//X0vFM5IYIqFFs8p4GNUno4Za4geGNBjdwHRrWQHWFMyXCs8l8liKfQ/TqvfoqKgZX
j13S2K0tb5+EJ/Ey+gUUbWkqATD/P+9M3Kd4ZETU7EqdvXejQByvKwnkckqTURp05sQADfogcATw
PnjSHBGzEoPA+AhLtl8AVpmH931NyxHrUZD1cpZjiuCPkzI07ENZJ+iCnjum+Suq90XOTAarmyz2
0mk6Q2RBTDVkObzeoVAK/NgmsqvqylYv+T0BC7bpu+At5+5dqJT+Z/N1cPfyl4va+gUlogPxzs/R
WoEo7HiQ09gqFQbSs4RmimlKvK/HFBh01c3zcCA/k5Eo3UtShfQYZBwNea5DRyIlRkWzJspx17Gz
EZi+JZ/JuyPSifDikfmQsLZwFpjfes+CYa722ryj42vbx1KQ1jDbCaY3UTHyGOaQUpjooYyDYb+5
45DTEdb1EBywwk3H4UCn3IOPmPugE+wvrehoWKvSLlSL2jncDOkNXJJEw6/ePvWZMEKbn9w4IXJE
VLNb3vsAtp7HnMbYxN0DoNfahKh1OR1icJZWwq07a9qrQbxd2bgm+N8vhU57GCh+LgjfIN/pcHDu
9X0BwUR4Yknky12LyM+pwFGvuTY5SR4dc6OolBqccWLoOYtZQo6AZyTzWksyxB8pY4MssNST0/Oy
ZGc3Tui6AbKYdiary45uLjT5XqovglD8rNloJIx4LaknxhGhtVCbQypmgJPgge8rPeoD2Fc3SlyO
3ZFKbwJSlFMFbrKflMlFgij2ABapMm/xwsF6yHSHJkWFeD5mptgu+gKVVNwQFTcA5W5/+lN4N6OI
gkLfJqcACSxOdIbwDKhKBGxce4YpR5ZZvIgbDXm6QG3CSLeGcBwXHq2AHNSxza95kkeTJKNuBPdO
k36YAeTTOpoQjjpNa+y48utGm0wD//tKlDjUsmoIppJn75Df92XmspplktC2+sjrvDWY5y0Kz+aa
6pkxHdlDdM1HNT8ophKx4ecmy5xhC219RbZR4uRzeLtCvzQ6MgxXC0m1znsxBWGqvHy3NOFQ88yL
eQDzFAJdPZTaE98CJWO3vzCK7cr9A1M7ITw3xGG2MfZ9f6nmKIPJ6YiJEB2zKpRNtUWwpoLtTZUF
QGQjWmEgjnOkkt3t5BSat7774lDaibXqQHrMOOTYMGXqBQIA4IT2i12QzBM2znkxkB9/nVBIiATo
q6k00U1yzEvVEUqskvb/84onuEQ5JgFs0MX8SC2FHddthWqva/UvIlWGBNxjoklmiNCctlhQQnZb
gPnRmDwHoGiq9FAjqetF2ebzzT6j7H3UvSus52cwPxCi6lWm8esD6TcUZtG5a5irSZx0ZpUTKJ9+
fLkfU83bQ4jCiC5eEi0w6AUiQaHqyt4yt4Vh9GYM4zTD3Mt/sU5gP9uMGfNDCpk/S/6cjkxBAErJ
gyEsIZ41+fH6zAlcfuM3rb8PWIGkxZ5rC9Zxzatlg/abNc6hUJ8rAhUwHLCv+RHqdisRdpeuYF2C
iPlYycnqxQxamX951NFkptnOAvOGKW7Qjtj4SG33JPoroUyLWztp+ajXAghyj0MUf+4LVMxYfUG/
19Keepknl5V7nNrsbqIayfEcLY+D5OKqKIQDv4t3qOhvjTQqi+UgDMEQ9y5rVCZIJIqb3I5VRSQT
0yzOr1VjvUtHbDS6SH/b4WyeVzwrtmEWcgdVVexalgMHj1Iikvtv5OA0m08eQCyQHVHiZLprhyYm
oQb3hh/O+Ov8oHQUJOiyY0GOpN19A0epU7iSDW6ttpvsEcsEKeVemiYqknJsN/2l8JrH6dZRpU1X
a+hXkkD/aK3Apf2iWBwn1pquSc6d1AYcWGRheVkvyBzfVvW1acctQ00ezgMTmi86Sfk0yp52imbQ
O0vhxey5eP+nuesAt9qYKpG2Ytoio6sbMVmG+ML4AKagbHp4QzY/W8QKdJKCV4c3a94hdcskzeDp
gX4mSl9H+mNRJUJfnexgJP0l+AwBYz5wQv18UHg04HNSm/j2ZOj5X3KGyCWWLohZoUZGAUG+kuLc
x1GX38TQons8EvmyCPPYXtsrCTGY/grFAindWOej4MMYjCU0fr1XNCCksVh2n05Y/EOLLxoPBGs6
50nwxJeYPfEdEoHfUQmWNF/EVKV6Z0TFbEox7IDC9MXiEAroHHGf2Lm0TAeQE6JmEewNw0Ev6xwB
zu3Gqlct99DcHzVgKd0+4htJu5Ey3tAFU++Y+swVmlPdOKG9CdjmkYBGv0x+E1MSFXYlU+ETvw5z
WkwxQqf3TTzYqHLCqtBi7mODBq4tVt5tRV/qQexsta3s0DK2PvExiPVuEM6VSBgnrsSzdqZEn0bn
a9qZ7merTyP26R2E0qQy93R3CCSf25pmTnZH3bBJjVnMeF8M1roI6orqTnNzcBFqVuTZAziD/cBa
AA4oI9tE2mLcfpWnmMRRfEjHwH1cCIM0GgjygfuBkWzni+tUoSYUmUbI43xZrv6QM06GqZtd2Avz
ES0tnGC3Al/1fkYojQVzrMbeRrr67U6U66E5S2dGRiVyfEDHK+J/RhOUY4ewmI1/f4qre+9+M+5Q
6AbpIaHeAmtQ2aQjM0VHimzDZ4gukG54Z1Y0Yblr61mN+pG5WYEtclvDCtb8u0+6WmolO7daQk3O
Yyhal3OJMG91XVJFstW+neS11pBf6UWhpeS7yVPo7Hh72hDjVeUu32tRuq2KfpPDyvena7QqRAS0
XePBuW8mnJoIiIOdPg/b/2dQTc2kqGa+qHukfLLy922NPoyXm2BQnTuTgmgYCjlMx1la8NH+Rls2
4oIf1smch5mfpQECPfYlh7oyoETN8JluK5RVlgXAsF6CXAhO561Xf2k6Am11ZY263Oceo8rNKARX
nU0OTnxt8eCCmaGc5PxTGi+Vy7nvVB8NPRe7PB8SWSmWDWr46aUF/fUoddGwm78dEsqlGSZvTR1m
v0xAFW6weRKG/rKnaamMWK9r10rXjMV2Z5y7aDqO42l3qlksHi7L7npaUABq6iumZw4CgAuBwJbY
oWtG2gu+eS6kWeW3zV/lSROiZV2P09dowA9I8HpeVg6DjzEEIDuU0u3gg5Ne7h14JU3j3loHEpGA
uANV107gF5v483TZri773EL215PtEDZbBirlziJvn82chnEnwBGKCUzmPr9toYJ5x7ovNk9dqtjm
whp6vxevAVxgmxX+QB4mNdDudPYUxebqnXojndt0kzvuBLP+NMPH0XPH8bjWGB1a5nhFEzLGEfds
C0teETgUoRx+bjznhRphSb1r4zB0dBbj5qePAo/1eu3mn1h/QDimQ+jXxEPMtbtR3IUbHTxDw7pk
TEzT/mhVCXBm639UED+KRJlBs6TJYSjshZNI1n0i1x6RkMaI4aZe9kKO/yL3p5nc/kHLhgsw7b5T
CcqRjZET+IAKFxP8+aP3Uv+lBOXQ4JxHrWE43DdzDHVoSCEo9QHvigtVnWrAzT19/lV8cytifG+h
yWgbmST6LnkF2PFuog06jI3GaY+uh4+j6F5FbDrAhBl0FTSOkP2UXdh8nwNE8SKy4+TZBF2xG3EO
ImJDCfZ5juD1MLEMvq+hsOV4iibsUYE+K8AePgWx2DAl2Zbj+baDKxH3x49nappD/gg48b/Txkeq
7CtG2JNtx25i5zuo0SZ5EpxesUNyUrC2Q5av05qH34ZQbB4+CxB/HT80f1pQJI5mHxNXlihDWBM6
svdIhZed5ziDXIddBwyT3LrQBd9D+hiaKxS34KDoyq4gZyGpQBszV8lNnalrXvsK6PO/ILAyBg2e
aduIfG1PZncCSff29QeqIO2tlBImx14hnmIjUMtHVe0jdYnutKgGBmFwLxo8xI5bvpE0zSDGRZ6N
sj8mlUhtziz/XXYgtFnQHgwJZFIPDvLSrWW/t/AzleTnrkSpFKcVL5dEx5AUOiTpbpT7fviXs5B6
heu2tH4TwZhlSp2szJ2Etnw2m/z0A4S7F60Fvkwm81REHXCoF6PwQbvjG2rsHgrSRCL0Z/OKk83+
oVBmA71jMLA3yvPNUDgY7DAimmdyuh7x+kC5BNgYp8fjdQYpecIRAT1EFO3A46XNSrd62op/dKVT
YWV1jg0vWG/VyT0PQEAhD8kGyDR5Rn6Z50fnDonRYwEn1cL3zMvTrcSlKLJIu5FyZbO+oGne+F2o
8BB2X2t4i54Fp/QFJ9udzcBrR26PmECCYz923kh2guzpgOAfKcAiJVtDz5AHtkFEnT7cBjheXk++
ojexQlcjdOVsR1X9TQekKDvjWb/lUsa+/Jutkp34wgbeNIIAABn3Dj2iRAChHVK5DrrNctW40PPY
05oXP+QAOiXd0/1a60CkeojXGLo1OLZxrGooqhop+pXPtiaobBr6Wx70zRV2NgvYU2YsOR9MjDtY
1rpcU4qiSGCp65R5Ng0SEVasiF6UtmcwfjVW59rToWlxJFP0BBCr7gtvvB6g2wuxayH1eBXk5HH7
3MkM9ycz8Mq9PWEe+zoWzu2vOb1Xs0bxtSGxYhVCXaolHJTPodz0WXWG4+juVZhzULNZYMZRSnb7
Ou8bYzP4LMrFAratnt7SZx6VTtDEmRfU3hkE3QBgqMEvMGX5gexj2owSjhMvIcrVK+66XYROGB+3
YouKPcbMtbHtmpNt8BRt4oLjcJRQ7Bk+S3PZnyNeK9UJ3+vCims8a8EIsXSwjoSGng2LGRVJyLqH
MeYoB5xwYamhXBa5z/OQoGxWyhslBnASX1tbL5qcCPuC550rzwyc8QpRggESNMVrcaeAwhnRnTof
8oplRs/7bsTkuR6KmQC6leOPGC+fhv74stYocWmxmVzHbKO+C5hDJEkYsPB2PwCq7JTWxV+z0AeP
/QLVzxr3TcnJmAGOLORdiJTZZbuj6kjxrBKI0Tm+r9IjsO0XqT1XZs8aa+G18oVcjmdsbMP7TeqX
4f/k13iwqlCE1Et1qhyBucGl0DTCfd7gd9q/2OVsYzM2ylWTwMeFzw+Ues8v9guHkvSt4SKWDyvv
aUepPV9JzeS7eEqYt5YxcwqLxhd+5lAjAxhmQckmdjEHLjWYZgSA5LkZYQkqagkS80+N1yvE1G6b
i0R/ZKKs42vifqVkzxAuC0nOSKMk9vCwKN8XE0Ie/J0F6MtCD/GYN05HsvfyTAfi57w9i/MdHDVH
MuamMQlYlIKqHuEzRHCe35AVskezhdu90X8M+Hh+04TZrzBJ7I0/OFh4a2Ni+V+hm7Mc8ayq2X7G
Es2bGZJBC8jss7jR5Xxqruj5px8qQavpeT1f6ZklB7hXjQuEalo29yG3BWdDik2K8rrSl1xdeer5
oPEFR+vWh0D6tK20DXb+OIevnWH4+XcDBbO1PXggN32Nyt+7H4Wr8LJ+vV/kxTlqUSolpTgTwKsm
Se9OofbsC8grNi1fNURg7pwJhnaYu+8sv5nB33IJUSwpTISK5nR/annbFD1sbG3ilTf/zPTHnzkk
HOoIwi7I5kd2lZwVMJeZW10dlOWzMxS6/DwAKVufpv6yh4QVhT1aoOBGaQYf6i1cDs3HdMaAzMEH
hZc6lyxQ/5n/268yAfVMt2knO++GPlf2INNKW31D+JmedPeQi11sRUoqZpLoAUrhq2fDel3tqg5j
NYksYSZZ2bGGrMCHPZ/Wd2zkVk69pL9oAPfaGJlYBQhw6ARJ7w8m8z+ElFgSm0rFW/ZnEA4qSAmE
yPicm3iKhmyP94/NYGFQB0yjU3KQJP6fOvu504hdRZIFot9wnrycDAOm1O3UEJGcFh5bjdFWGbVb
MbotcCblLfv904nf66j34Y/STvOAyUlIz98SjhPZU1ddoGJ+/KmXZ57f8Wv5iGaY3s3npXBanp6y
Qb7S7HuNlWOCZWNmIzLdV4rzj/5rwaXXUN7fLK/BUQ3fkmWyXLbRTU81waJn6QcbEKUshNC3iKuX
IrFRIznC6g4z9YKfHsjCxayaM1bYKRo4sRLS3e7ZlMOPTxB6ndOYx4l1lZOCFkGovzNbbDf9H9Dy
TxX5jmHtvGg9u+DPDqmde+p8ko8u02eFMB3vumLtcnGraaT/OVmjv7xUeT4Mzd8X+DfatBFeDArM
Ddba5cppiUDA48h/vzleJ7NgBAKTlKiJxaVocwb4KVqH/101l5iPY5GALUfCW1LbgBozZWaMAF55
uQ9Hw2Pi6q01S3wVsMCU/QiiW4kd982MoAPopNO8gjH6gAhKWcb6xYtUR9kyhOzu7JvGKftsbL3u
djJw6EMKN+vZcHgph1lAmCGe3OBbQ04y25q4s6/H6mhF5ka+t7kvOzpsDub7mzQKerXY/a1MBjv4
DrEXpzGxu5tULmyaUsAF6V20/ZcuQcurbVtD86oYY8zd/vLpJhDgiE07K33t8CGKW+2aGPZLFPTn
PdfOSFf4I8LIJ1JFb+BMvZg8cTUXUTk6AHZkan6Jikj8dES2Ft1RJqOiWbyWtbmt8TrpY9YrqAY0
Jc6A7gLPSGvaH+cVECKujN3L9fp/os7yE5Mfr/ZCBOZFsMHeY7LVokmhRvIMlkAFGrNgSgAVVpkj
DfxtQavqkGi5URjTyVockj5/pAf/lCFGyrvolq/ry1+QwPsaQgi6aEBz7AzxIi3T3PgLa9Uk6cXy
4Z7MT8IweVPBx3GqU454vCAqXaKe/luF8c9u2xTr8RwRR2MYBZwKQa9iUT4QESMqgWE7m0LU/SaL
aJAdvLW2MmoDs+ulyGq8ZAhQNRSgHJNdW0RR+Ft8sFp1ebUL1LOTs7UHkjL5mbRN2jtqRORdWXk6
sZvC1UUgm/VLio4il+rB+qJpbc1AyLYnrEQy7KkAZ7tbNIJB9VYO+YQlfmr3bzTwymMJyw9gW/wz
lZ9hlLrpwN+sQk18FKMb6KrRsGBCS7pjht/fjmsocKWJmoMbdmoCRbpwMJqBN9HsLjXxfh4YIEa7
utmtNXm1LG9Gi4pNDuEubSyqSRf//nj8pOZnGl15eiC01VgCYYtUDUe8fd+fFVLqHRQOiiELJOZN
5jcgDDC+c9gBfQ7rS7j+i9di9gDeMS+r6Fg4ijuvPDHZX34KILgyjlO1kOvnWY9jC5VCZouHhfa7
R2yGEAMGqC9kOCH3G1lSqGodh4obkfQEi/ZRM9dYorXS/RrFoECIoI6cuR7jSP5qKH32rk7z6DBr
lloay5+CbXCHYMJJnkOgab0DegWRoa8URDvKjK3wWVtQjKT+gXq50z7rLITJNHLqR0OTZ7dPgBy6
4sP3OlkOWe/nMX12/Ja8Pf5iVlSFqmlq3wEDg0qZVxLGB0eHzJ1KXRVVN2uGcL57tALLKNNYxMH9
WiX/862YPAhhNpNNQLgDHLeqBDGcPoKYE3y+6090Iy1JirP98NJIaJ42tVoQTIy2F/ooUMPGD7IV
trFVy43T3VJCXkwZ5wFs9du6csxrVsEcqzHh1SvhYp979kXUWis/eV2MCdAE3DdrexExzQgAB886
ztFVMl8DdP+mSUvqVZnhyyBnwxgp0K/z4w6srNAnrCxZ7tUS8/bJWlaVkUv1j93eeNgptxHcmfPx
yiB0IbutnIg6cMjYM0ggWK93sxYC/Um8VHg7oNgLRI9pcKZe2WQT+KF50jV89e1aGmwS18ZIWIiS
0dJJ1jNNDylCzH1yG+OYUNPLTGn0bBuqEo1GCFx5SROwz4RXsY9bvWvY8nIyXi7RAguqzUyjP/xQ
hPmQlZykE7dkbtItqfP1r5cYNWcvcHBS4nIAEoppPOsuTP+aVZLSqJc8/aErWVbo8E9EYEyid9Rl
3FQr7WauafV92/a7mcZUSo+1rKJS9mDGSslyzPKzOgjITTlsYjWk65yszB8agDiUos1wz+feemqo
4BeSx/S8O5YUS3o0EMBUjwtrM4CH+ub6ZqiYRDvUlVWBT4bsrJBAaWztKW320O1a9cFTMB7eD+ix
esG+MwCewTu9hCj5MNZN6CS7Cn9DR2+721P2nB7mJGqQitsjaqR+IRQ7JGHSFDG+hqzxM7S0gP8n
u79v1I60CElgsvCzW8hv76tJH2PBqtRg/cPJ2OxrU/PM90XFQtE868U2Zf45bjRwRFzmlO37Gov5
w7G2ee0k9eb0K57eZx/MpfO9hhRa0ohwYgHeJ+s602YBp32lNVF8Lz9bsRTJHa+YGI7w6c1dmfcP
8aMvdedpIr8HSLkcvF7T85H3RuVns27oF/e1Z3/qV1E03wmYjDVZZ9LbuFRmsmhqn6sJV4DpU6mw
0MHgdQpZDibHoxGoXKYj5nPMwOgUl/XzxnI4XeFTbRJTJ4pGGmtoJBRkxy+Q2lawZ5LQouh2fkrL
9GRG4/CTU51pAirjKChA4Zj2AbmfzXm65lyGUdXLnmlRg00wtonJP2QZykHURAHun0M8H3/93l9N
OehnrogiGmeoxNp86CUxhPOdliT0lqtuGvYslEQQWfbBDYO3+LmRRtT+VRsCZZ9byIy11CtcrmVX
lw2oMLWOJiTGPBwo/IfbekJW/a2O0z/bplYRN9ubkNBSAQe/vCv+Yu1883N7Zdk2jSMXXS2K8lh+
Fs1zudGx0Lsnpk2EwfYCOWlxWoKN1PDk9xE2glZXsZh04lbm/EBuhoJSLxjF154unosjpjg2N3eC
AWDOKqMh5M1irJvDWSqvk24ab7B9D+XXf2bxD/eTinfVEGcB5edbWemP5EDjEG5ij7C1YSwKiY4x
tfjZETaaSRVEA5rtXm2XABVX57wHWL1tDGFTfohp2L5PXRSTjmskZvYzsz/5eDQyJaFDlR0wA6NY
I6p66nUPm/ffjlAgPasioVnFk57X442VcMg83unY9+ajkvnh0aW8mcRUDZcZGU/EKD4sHasvbcD4
w6nyHE6lFfgYM/jmUVQjX6NHMvfBMROl/k217BOdaDM7F/ylOPHF0FCLwt+xjMExoNW29oHlJKDZ
uHv+vRdRD/UYRASWlNzEf8gXFXXX0m6gMvfulVA0cpQajj+ETkc+rqKAsZ7WPprw7r7bevpAg/CU
0swnbpH0F73HDYDgw+vJGYYP9R2rXCEfW0JaHqRKUiT6W9adY1GqEbS4SVK5ESuBZWkzgv0Lmltk
XRwpXyPalDch3Wf5xJ7LCkIwS8+69sqdpSAcYqbk2svE5ydrhVcohrTs+8PqwKKaptau8uT3IrDa
ev6TYVRFG7saP+HfUY2dRdLYidRzkiwX6B8Hih5RDEAo+kc6ndLZ2EGowP6yfCLr8t8yOLkF4nv2
3/tkcR+i5yliW7CE8/KdMAyCZfyiqwYIHEW5ZsFa+HPkoF0l8TUG5HfN+ppTuXufObMFUX552YSk
4fqefbLHGox3ksIcBmCAdxnbvT6dt7vvBxzJYU/pMo7bR6z9VHhz8OQahgRUhEzU1FfZMDlUgLGB
pn3O8LltTi29uzOgR7TWAvkOIkoyjHqaKmTZ/xkbeTr/gA/zZSFc8fGCrHkZGikRDL4h/L6BBwj8
BuGzJXbpPsQ+Ae5uYS17oxbnrwZsHtUwSiZO+42SA3tyyBWoYu+MA3VPVFlwQOLHI16GNTvSldVU
mIhWX+jLYTigd+gyGHjYd3+A1cS2vPsmnN6FG8tgvZF2ghaJRuoToW7N3NIfyWXx8TtVEorAPXSo
WHyFaob74ZWce92GuEquUHdG0h3Jaco4BVSq5yN+GFHMTLDQXHsnm8JkctSqPb4Mrkju1qfHYkXM
y1EJ7LJy7oF135aA0xusgR1gEEqa1LyWgBkHONJ1Kc3QS8+nvdEdX5pGD4XuioWI7jaSW0XdLSGz
3YbpOUlDZ7V8StzDIFZLF+vGtn8CPcItdBKLnEc8be8JvKWXfMWON1SJNu32P+K3jBLsZzydDNoU
ym1pGSvblrldNuIqlpkCeyF7dQoaOMfnNW/qDhJiKq2dKhpQl7WLbD9G8QTkcr+UQmj0G1aNmeqy
kONHPXWG1PE+wlmTUJKx/Q9nVM6pIOP9YWUdpYXbLv4or5MJ4gmngiaxhBwPwVZtDlTXObKVEqKV
NGqvCgZXr/wToVEraz3cLT8WfIXYKOplycaIIneWkWfMyI6fgiUSUL1o0/zJoY2vbsxuy+tiWPJd
+PUPmgEPd3DqDoEChlDwGLdKwfUmzKPVbWGzFKde1pVGEv8Ek4oPEk1p/Zvl8MbeaLvCRpahvzkH
or44M47AgZ8pUONKT9+nn3Xz8w9JhvT7uRtnmfY+hiNmddPMRlRvtgUbP2aWkB+ib2/0pN7Lpazs
df06aIHOuQ/Sc8hQkphbDh5N3MBVX8SPftCVTCoNJY33bdMWXyMZHyEQ5DD8u5KX8NTgomj49yhO
eJW490L+Qua6+i6yOmMjN6o5HFlKLMfb+ikmawpfcJs/8XECRuZPVTy7R+invkXEPkJoET0cTAi2
vub9lEwsjjOaEd8eFuprQtt00yokJ9y2T45ElXXcFsPyFJnNJU0idNTJ8mk9/azfy/12yP7F/rKi
bIWn3doIC9vFzqAiruLfxoTCOIuRPt+OYir5opwWGEM0NAu7KQr3AZPVVMznhzoiMNIa9CmhRikh
zU6xvq2eazJ0GOwr4wrubueGAAteDhXea+ovGvEgrRuFWho2iw5cWFULNLn/u/ycZDS2Wxlqo2Y/
AyYRjg1Ay1SEPMPb923V/b6r/Qzvx9A71prJGB2s2TOC+s1jT+Un8jYyH/V26Ee/0GwdfJwRybBw
/PS+1CjgXzDPOJxa/2ErlUQi/oT0kX1UgrFjR1uwfSMmvRn2GOsnQK7h4b6QD0z9luxBKAiOgW8w
Poor29qO0A+5epLd3CCrbA8DQOjmZAvyXb0+Oy+s8qUTDcjB1EIE4R+9ixOAN1hYXGmVoy8JcpCK
Omj2zaXOttfxo5U5K8UkHYVhsGDqp6waynnC/VTWmpRtVGY7RJOtrZ4JJ0FwBCvbooocoQ/9k7RE
OF4xBRMbVtvJsGh5jVmdo+bod7/wmHmtBBrEH2HM7LkEyWCRu1Sihz54ozShHyQhguqQYp1voTX9
sdOCDhPiS7DYUDFc8OpTVCCbms2YztbbclDROdygfeP+AV6UmdF2Z8La+Zzh3pOkaz7Z9Q5QISFE
gZR8HpJDUQ61DNJvnBlA7h9RxYj9Hn470qinYsxf1GuyYmIHrGSfKo5G08dIxXzdp/fM/qHTfSDo
ePSAyD6+l3zrfejfTicTWnGNEu1Lc0jgrG0pof4VDwDf2JEAg4fhJW8CILq8TklQim4gTBsIKtk9
IhqlS8FDBXvLlePYy6n8Wupa5GTg2FZNr8NCA4C4tp6CxJhf6VKYWwP4+y/0erBrVy7YnU5xkdPY
qoLNKhp8QPvV7/oZB0ZsWT7wfTcO5eV3hQ5/TOqSMX8ddZiXqNaF4GPyKOCmF3i8c7befAaezT1H
Db33UhYxFhjeSS+aa1MQCWEsoCaiG4yoOKZhcKEWm0BHSq4V0IHALE7MPV3EPexHupcLCHw7JFgD
ItYsPf1ZNBt+ZilIyeHwy82NOyikQLtOwmR2QHkoK4ZRJ1SA6UO8rksS1ro9g0/NIRkoINJK8oFR
uEdIc7MqjmrlQSqRKTS7DEInPzcs2mbCpfOUj+QVoZbPWtLHNSuqKjpJjZmWOcPM+a+71dRevG4a
erSG7dS43s6Bk2OWicnrzFF0uFCRdCt3kaoB+iexxDs6l9D0x5iYk696s95JiLxkyhpLIAHL3uP4
eIzafgVUyI2Hxb2wgLbAAiW2es7zcNUU3kZlHNEfGornrhnfdAj/N/+/ogB+joCPLJR8v4M3Fw6s
tNuz9532uCeKtTBJgbyzEkSYZpGpkhzRXbWDaGamWlBAGKcXpEzi5tfHJ82gtWA+gxnxzWfpvBlG
Zxb6RGCI4C/EiYS5zqWKdcxYLPeWBSiqU/6DVTvkvw4J5i9OgVeGjU5y5NmJaRKUChQpprmRuW06
R0xGM1n2G4oakXvdZuz7QjtDvKZ15Dy6PGTPeqFVariMaJXlHeHmeguurlIZFpIL8ZQ388WK0eRR
GrzWSetSZ2CWbRCtTyLXaeRLt8GLS+bnXTwpKIkps4cs4jBsSOfudmd7RuwYOuY4A5IYB72IShty
XLsPCCCK5KyCVNnY71o6KSNBD7IVdb/PY+njFJO/de3A5U/32NfCwi50aKxXigIrfAD9q5wSeD8i
vaOgSYoCBSjVHo0Z/jzcgDcfAayCoplbj90/zxHHjjUQ3dZvUVuq/S9yVVRn1yMEU18yOJFgpitc
LLv2US9PgLMXCkKGCwV9KtaVSI7soFRX43zcSqDi/o+Z1ps1cIIdh5cvG5wD1vguiDaLUBOFxsZI
1IPsPwoQlvFA3Gc773ivw2wJJfkyBbTPlSq4WEDYs4mPlcnseQwrp3K8S3CHdnoD8ffQYmChpzc3
NB0sJi8jCa/UvRMiiFEM1TMPiSQnB46tT9cIUktNwo9/rAi1RW6B3sbTSH4T4BXtLJzkB29CibIf
rtRaVw1Sba+W08aXmDxFzS1rNsrp/NfhseZmH3UNZpvqJSF3XSYqVe3madbqr2eDFZzJw5YiSuzd
hkuNZL5L1GTb0dy/luY3dDUAafpKgXY1xL2CXov7JIKt67UxS3RZqBSn4aX4QyLiT2JrqMbQqCuY
K28fQckGYu18s24MbJMv6MAPKo4MiqEhmNruL6DbMXS+RPrJvAW2MRlSj+bBhqpiLWjq8z4UkXTG
RKNOlFUbIkjs5y05goMYM79kkMba1XFDY5bWpSPk2BCikiXS28IoiCqLFHvhqavXL9ikL/RXv32z
nkOd/68TWx+mPYZarikNdh0S4mUDJou9dNghFBCcCEjq6jdwZFuR8uph2b/yWkFy/Z649Bjk1kZ7
uNNaYegD7eRzqychdUQ8hpj0Mlkcwx0DFh8V1buTFvxqcIHrhC2AsmeqUZdwplUucr27H9Xmu2y0
tejB5YZ3A0VmR+3qSWbv1dGF3KDozOitWrla51JpHS5h7t1Wr/l7/q+MjXzO2LDyOL+WAdFCt8ft
g6oRLwTzYnf8gjAkzkEhwOQ89iENI0PYmvh+Yeh2U8yRQ0TrL6jRS/iiR/WZCUbAYdflph8coFkB
Mf/OHUr1DvF0aGKkWmzO6r349SL+eOoMZeWzyqMET67cma4WYqRC5Tp5QNFHTAQ25JP8V+/7zsC1
XK05oz8giggV1364XXNcG6JsS4pVrcRfuI3t5SjrKkC3kxKlOyUbTdBcxvaUb/iLegC5rc3tUi6E
NJHCnGM7cORLBaxB/Zy6O5YEmXoWogSFbQW8KlsHYB/diTEraqBwdPci3L50Gq70ZR4jmrhGtl3x
7BM0tGWZEJSuZP59UJrJ3ugVwkyuO8vQALest1wvMqdXlvrssuh6vEUgUElEqXUAaV5YO4AFyvTR
mxnNPWjZc73829KWKqFnJtsZdlz+gf9POu0e9BxEZh2B6aMEr9Drstoo5dAMmxWEMgIKoiP4gBib
+Yz730GY8qWvnott9ahDqzMlmIIF0PFRmXnBNu3hz7g9GApTjW0XmlSegw3uKp/8ATAh6Nq/bkB2
Rm7PX6h5UUo4ig6gk2GQGokpoLptlA1YsXHlUGsEEOEwJ1hNCTMdBYl/fXCXySmNpLr3FLzEmJm6
6lV+HGCUgMTDCD2iV4PukbR3+qGNud5RG6/kDRuHORnxD50dPMI33q8rPqQVPHD4KvNjwJmmhRJk
t6+6ck/DmpMxYCOQk9GyWOc4s/x75b5Z9dz5LZScQWahsYKqsJlwb62hTvtK21bBboxnWZnTDRKd
Kbyqt3s7FL8PObZUrjBoiPuloTPu37ZwTGxpJa2Sb9fR4ymgnjvN8RXSY4hV0+ojndPl5u/h5L2c
BX7BE4jYaTHLMploBHAYpVzC8wfkOA0dbJb2//ezerIXZyP7680rDiDp7iCpuFmrbUl62Xx7Ww6f
N4JIHLyGV+xobvQZxEVoN1FGXJMokNGjz35Hdfzo7PU8vxZjSGamNhdmRk3GghTmHZjSYKQ4zcXm
lkKDLgAf3KGx2FNKifDEmQNIZkzDdmuKUf9veKaNAXpNpk9vzwO6Daf2d4fC6zAUC5IQP/Q+Ba9N
6mcRI+8D5Ay6728fYST7CWZbLNU5EdO7/iGwTRQNEpvk1xbvTdxQTWbIdrB1LKm3/Su2I7Fn1aCa
SrOWs9j/RD8VWzrb4iAz3trhy3VJNGaV5sW9yfPkBM2rnrttyb6KW8ouJ90tX/lUm8WGolcEULNn
H7ENRJ9I2DFXsTy9yztZJNF6lsP80IVcUk3nGlKpM7IGBnhgqZQ+LWJQmjuW/WxHb0CXMaxsxn3F
kPDX/DH4m8TqBYE0hCIKvgZiAW/gJ3dm7jte+5ATEopszHg2o+3DPF0MR0xhsWMroBjDaCEv7cB+
fGgA5NelIaWR5s86QpFyXduVySM9uwgk6avLzlRWpNsF8b8SEYztCFms9YNq01apR9Tl+w08JD9j
n1wMfPZfAGNbtDQfG4vSQ7DMX2MxDZ3oRFU2c0iFPoiJBVvn9q890AgMMn2ihwB8MONBGCPYaGLt
8GuRP7dneXYiXgXkNXo11WTHqaTzbqmWIkZnYvGFXP0VWFLhzkut6Wc8xLxZBQC0q5ixw1OyNojO
ryFi52O9LJ6ph2ciOJP786mFeyAHDAcUb80ziu89ZN3vfiBaIR+M4L9YhnhcwmHxoQCekV7Qvtqs
URPQYYSUXg0fOYjWYB5bnjGtU5lVbxLZIkfV13wAyiwtfAs8iXiPEFzr6g/iLN1hfBZKXRx6g6lj
Y0aueQ5f+rfGKnRKyeXoartkCJIIaP/ueTDCrlP3/SjRGCPO0q4IDXMdWNk5baR0rLKWCB5hjfKQ
gp0ovwRvXWm8cs6r8gcoVFw5xdkAzHuWkZIDKA/tHIq7mexBhPWBD76j3uJH3ltVYxGf4tBNyZj2
FCyF3WcEpNpaMhzGj49EhTnnjKkXrqaoJEZ8RlHOHmNTQRrEN8ODWLfy65Q93t7Xnb6E2lGI5BAk
JrOLeJXFZv3J3GK+3O7DQsQMxz+mtICTAuD9tRaSYSZQPGcI6E0Z4P6WeWktNzeMzC/5H/JPR0e6
VDbIgNuaeFTsWOSZIZM2ZAElPCjK7sfoSaKdjbZOEOdzkdxLMlajgUDob8doin22YghdFGF1tlDa
O4wdjnhJ6QMbmn+e/IFinyNdv3fQLHZleMTSOsGIm1E3R4RQR0BGbWqHkrV2AX7L63w6vkBKaftH
Mu+YOdYf2hqOWtvsSyGnNpLZtEDhTMSvygIxN2NlMpAjsMzgmNSNjuL4KgUzdCFivTmqdNYtEtTV
cOCKFXlAYFwvinPYTgcaUgHMAzzqomrdbwJlnlBnfu2ZjIeMzc811vxdSbnc7nb+7zigN3e9Qz+L
mzGQteobs2QcLwtH22m8hNHLgeY8PMi4zstiknh7LIYOsOT2wzrp847FyAYnn5GJTCky5/m/IPqG
E0ksnfp8Lm69WwBB6pFcvcJt0IBTprsOFzBdZQBskmUq8GnoyEIhkMY2Qj8HVn2IV+DxQhKNLINq
3AcmWtV7w6WYO5ciFRuXWj4MHDGgArtpYjsndCAxsD0rrDSuvTMmaW8WkH5yMU/3PMekQlV3NGCm
cXoxasESQfPrmtTm+Gt/gM655Fqm2hgFFBlBDjlWcqnRDtlpw4RGHZFgUBVQfqgqS51G3bBgULNf
EwFjBPO7/Mdags8I4/zChCtIuGpDpAyNzYHo17SsE32419LeP3LVN3bdTjRSO3tuZaQB+tMlKyoF
633QOIV1RLIjRGQk5QmIyhxQm+NQua2jlGOaZVJWVdw2/GFDGsN757/JGEa0NAMbE7EHrLaKbyAx
U/W1xF7yn9tQBqqzr1K1huLT4SZYq/fi3nb8CVypXBtlGIvjtg8MneG6bwD7gSEUhDqZNT0mQuVq
dawMGnYj1I/3OiiNoOWpsHogL/LC+z9lMuEwO/LeBVGF0MaVa9yAk6FS4wEE2W9E4lFFwrzeOVpB
KuvVF7xLqwVc1ybjCMcvNPZI31qP8yhbH9qQO5y4qYSEYzZmkDb2Tts/iiAcfB2CoRBMiulpL2tp
FQbIBfXRBDa0pSH/m5v3p5VQEH2ugNk3qgh56ZF9V3c2/qvhM8MnoZ9FNaPdEdNTakD2pdwNt16U
wcqaT+s/hgsKBjOLTyCIuHLmZL1en2sALITur+b5WFwYrZIoRAT0nBON3rdpIKGen5Q3e3+JbLQV
sEhOUR5Soq+Po5aU6ftNuxuTnq1epDZjB5Y6PcbSUhE4Y1zYU8P1Yy3OvSFFinQFDc1kOr43aYJT
MGc4IckUdo9etp4a2gROowzK71qVEP8NUx2AToMtaXYXulW4Mc4zgp0IO5ZOppUUA20o0artdT8Q
XMDvd16FEotkq4uSxuHHCwBTdq6DCRTudrRXqSP5f6YjwEKwg59UHBmBj2dsadJVoTXKG4knfQ67
QX791yI9BT7k6cZg1YkFEdL0dX4jay7LTTE25Bq6wvI3XPgH4TMOEnjygFbUcWAqrHvEOvaThCsi
Q8/4lnV6I9wRKUgauEZkjPBjOzI1W3QvfgVDu3sQKTGHrgAFcqPD7QMypRr+Vsu5evCwjFcKRij9
TZRh93/AV6V2B9sX10EGlw2HXiOnR3l6FUaSF5kU1nn08rn2SJ24GxH8xBbQ69SOwpTdy3mE2AH5
Tgosaxdzjzl26UcZj+IvXZ9WtgxRv6kHpkMMm7Afz6XkXm2L4V18YRbSX7tHjvFz3OFd2DjZy7Zg
ohR/IaXxfrtz+OH4OGhwoJNZ86vaXFxspabswENR8+WSbNDGqIsofv3xobwNoRUBZht/TqbVhoqd
MIIenShfT8sgwKN2Z2k9NaUvjpLloOx2K5jm7uU5opuPNbmU7Z7yKvX18/9U0BlxBZQ+fNhMtcDQ
G3pcyIwlogzcUbcg1yaNTB6H34SpSif4VZ1QVbPGhb26ax0tEr+VO88KfJx+2Qztr8Z0LkLho7tW
OIrIqWNRZTeQ8giGlECc8OiSZ72OrEStHh0RMsgQsTEEr+zIvuBEEZi4vSgYEbqA2g84gOAJmbIi
t7Khw3sgakVtipPgOH0Zi2iO2GUzCzmnVJ10S1AnlPGF1DopUgyYTibh75wHpzaEiis6bCrBIlD0
vd3J2n18BiZp0OIh9jChbCxvcTRVe/W9uLlWZx7tJNd8QVNqWAFgV8Kcn4X+BReaPElO7vSsW95A
hAXPYzqve1dgMRMGSSsGA7n1Rdjvkj7PTYwSfBD7fZf9P7FGoqYEnTdSwNT2Righl74QFDdrvK7n
nnu3bHb1MPUhzwYsyWzfMfEZU1XTf/NINuQipLW6rm730F4vHQAMlW9f5Y3iYQZYJ5KfU3fYvh9m
VDWvwFBHx0Eb9fIFt80rfbHnQUuiKWCU4LhsMkpIhDaqOmwjuXQsUUWTkrf+rGhEjjKXedEBSNKq
66RunzqpXiLToZkwiJFmSs1Ntol7xpyvcyDWYjk/FrtXVmjxSG4zXdPknc+FeMN+rVzt84RMJmpW
JYpFIOtaEEp6heDOFvsZ82WDgt1FDjj1KcxmgRcS+Biney0tRvvy3xzNgP9SLpn6ZqYnPH7Js1kf
MWvrWolLAadhnZuMfz8EscRM+26Q+5YMxUAD9NZsZK4hSnqlM/D/KKtaB/8CmLZR2ApMvFHQDFKm
VJRNSayiwsTx7hSF1kIYYbkmUEZyyAmT4ZH3LGeXQwJFGi75ZbT0HEiSKUl4ilmW4GBfTAVyA4dl
t4o8ict9UHXbSUsHPsl554JDDhE9DgTF1UlmZhJvWc1rb1l0PMX+poxjnCbn78umyst91f5TsU9Y
UKzbaJyDvrqwrSeiOcECcNq9asB68rJjsi5CmNEgmIr5tNhfKxYD4pdtP5nMRY0FdQsU+LVyCrNh
VFun36lQCOQF7RK4P49P96KT8NB6w7m5Td73I1ijeuN4p29KvS1hoS6G3gF4qww4cTGBJlpjCZiJ
ODAW3HcRczigQohLdDJlIOkHoXyCoSx4r+IqG2Nod5antsXG1WEvJdseWpsbhFjudi0cp7BGLCpL
xKocU6Bckn4y3i3nQ4dOHZYc16Tf2+WGRcum1Kg2TyOQEIzlz4kz3MvGK14hLaL81rPJFON+OjWu
oBCEuABeo6LANQ1SnzvMxX0nyYAN48UIwDpx0VPStLmbre2Zb+03PGlEFfEMmASbyamOm+/JINhD
ApB8qmHANy/0f3HNalji3MEblvlHd4FwsTOImEgOunIAw4XmpPC6V3o5y20siIesXbiY/hFH72TP
vjbp3LrUj8qbVj34HW+QM0VJyvxaccj8EUdxQ8vsfF+p7q/6/M7MLkqVBgJY7csSHMVftOt2u1E7
RDrHzfvHfnVKzx8r6xGt5Zz+ah99sxWknPWDVV9QXPm0V5qHnaIpYfew0xaiBcnUk9P6NPZvvOJ2
DSAh+7kVEQGDY6lSuvw0FGVD6qFnZeq/eKzGJRwrwvlGQ0hBiBnGSpYc4Q4UoMSQVMVeYSTz+sna
aZtrMG9GU4jDmz5lGGW5LdYK3FxHn/m8EEKkfS4H3wyRKCQh3mboAImf7ev6aObfnqm4BzUdvHS9
tYuB8bCnpcpKGwRA0d98IyxF+2xBYUGHHF2V3F21y889TSMODYJKeXA70K4b/fi2+PckPjXNgpFJ
cIe4O2yLpifAMbt88Tbzw20ne6kakLY20FjjMWHcAwaJjkhpJlOSdjGwE0+USZKggX8CvyY2sM/U
F4pLoUiNpp5FtFEBmrPW+aUtFtgDDn76i+71TOvmCR/KtYjAcvPjvaqAmmtz6YdgjOHXurbrXeR4
xfp68UOEgEpYLLPWVN+lZpPwn7Y1kRF8q5Q6pQe2DEFBAO/r0CjeBW2yUIlPN0HuamYzb/u4XAyg
Xq3bLVu2NF7I8vJEOSZ4LCNPLDAKXKKoukr2M7/qjnlG9oEAws3GCQGkSH78XEQaXvflAUpes6C2
NDlMYhrUl0RToTSTAyklwtf6dLlCTl4KNXP1n5x1wO8xt4gzhSFzySvKfMw+/hKnGcT5vsYnHzb0
B2ZSr5PW0VZfmzfeBQ5e7feDZEfMWEPAEfG9wCPdhFcSbqeoz2u6FcPZsuTN0Vn1lvu/X0JySRAC
C3i3CJSbBoYnWwGw1mktDKlRvWQ3V+k1ixG5WPK2LKCZKZ2ppEt2q5Ga2FDTph3+QectHA4IvpMp
WnhA2is0JcAHqrIuluVfPL95eHkxM4s6J06MWrPT8RMxjlUH/pGUDRogT2RrwyGINIJCdTLJx5xV
u9/skqWGg3UZm3qBx2+En5BTTDl1tQMjq3meX4vMU7/ZHw6sK9g6uKsnjUeJj8VPUfmmri2mDcBq
+Brv4TzxTMcvX8OpziuBP8sW7nruqArTfCi7e4B8NW9r924xW/OybhK5HgxkLuf8zx49LtR4ACft
pwrgY2wWj3Usgslz2OliNiN8F0CWErDLUlZTLbRD5/qrXJVULXwOF95uE7PDEcM36HQsOcE2Q3I6
aJkFN0AgtaHOie177AFWr2MQXk+gXSXeucHa7NwJa+8gCTBK7ZPLmgAaUv8Tr7a6zfTXXO+AzKgb
P4e4AgIG+ND7MNJQhAzVweDHCRgN8QhV/DAH51J6YkOwEgBtIQK0AzTQtftc25Js8kDj+GKLJDU9
Tib6NzuXk0zq0UBsH44pU7wBEaTGkDmY8tlcQ4yD4w/vVwn3BhbVT71LB+/JybIIGE2uQm58UHbW
QHLDYO/H5c3IMWnATrHJ7Kma2RUawbH0VRQU4P7AVaFHJyx8MQFBY/VnVyJKboKPsQ5YTzvkEiTT
BWY3w9ew7ZWou0hTUKUT5K4FIWOCxi9O9RDQVDQuHIqGeJQe7ynaOmr9jJiKJtGUOfsWuAGkrV3w
0FBCXjY1Fi7UD/hjwrSKQ3PwNKcjGO4i82aYvDIKXmCAlDbkw56woLmuPqRcuJnvJQ4mLgy8aBeK
lLgSDnNF4/osok0P7/ajnJgA7U6rCA7LCcJqP3W8qyHEWvfvLudVD4th+ULzNlQpuRQChNQypoWC
WlMqifOz+Mxbv11JFFVnTLf191rMR7Ble1lkVta171wuc/jrHukX2oWGUHZ1FIgCM7vpyGmh4UhC
kn8cb+BkK8hTTC8jTZBRs2tl19gf9axBl9pMaBkhlIKn54rdxYbphbOpZRY9XdmzKbOPVL7R7Z4h
tsawg6OK5i5Mmud6kJClQ9Ca16PEVGAajbLzCk0zQCKhZgYV5BLK/bktPV4Zatz3Ji1OpC8u4bW3
6cLNHADXXlrHEAgi/gjTpRWUly3Dp2VaC5Bi1rM521zfaYmaOcD3uJD7+DvE65MLtgD6GIJ00LQd
ZCoXxl5zjkgjOTbHaqrG2NCuTUEkImXeAfxGMw2lueQAKJ78fjX5GJPbUgZucyY24q13RtDHpx/J
JlfdR1fg1ptuKhTTFVshy7GKE4ZYzNn0dQIukEnSZ+haPqmDhMUjVJTmUOyqnTSJzFxBW1iXalGk
MS8oxdjdpuAq1EkrgFTq5qBH7xRIfl6w8ZtSU64fmZPw3mHKBHYEyeYhZaHJ0N2ZvV+AFgigw8Hz
dpq2qVJDndLZ4ndl76pk0oySicJBSiv/BfG7Q2y2DlQn/1VVojW9ZL3U9S2xmltbBretl47pgXM3
TdPKPJE6ny01LVb1Ws1uDMHKnynRBAj0GoZOnVoLVTHS32Mz3HcsxfH/kTM1Sss+pgtM3UfZ2piT
CkWndiZGS/HgaaOAvD4CDSsBXxz3doOjA3oNrA+6R1xk2uCTfEgNMY5wWdB5Ou1Dd/7gKySYeFqq
w9slF27Z7t7dcD3WHitJO71UGWlB7Djz170mK6rBZof4XC+UBDl3elr4pYGgVKD3kivsZ2K16tCk
V0ni/BBputOmDIWjCoCntbF+Q0lZAdCrlOFj3Jc6u1EzQcHeCzpgb2qlws964WDj/cQUwwUdZTX3
6rjUcNju2mKBADKHOL9TXyVqPxbfzeu8Itwto2eyFgnngk1YX/5x0oWByWwcZd5PW6RUZrCvb/dL
nDcd/oaWmDk0J4j6rGsFk5JjW/qBI35+hAEENPbO4RvakvSJJ7i/igrbEE+wG/iCnK+FBgnrgbZr
mIm09LwHNnWdgoLBgMNUBebhHzb0+TpxB4D//ev1dLSxnFEOThdJ5da4Ysg9thByA+aJx1elLVSw
rNWTFnPuyOGhb2TNlh5G8Guz6SQCOZ/ZDqqqmwawn6nX+LPpNkzeoYpEhmsWBQoZWsDONQwHBtqg
/Ru1E2YbHe3cFhGdfvJyNI6DIL7foxcm74jrdHvFTU82NGmKADz6feAl650tpcaRX2cuy/vd4q2z
zGrA1VJl8tzjq8WuC8nQ9ecXJq3ampuMdt3X0FAqkXJq/z5ZZjo9UqW+sre4iUC19sjCvRiYSZcd
4p0zZTGX3L8aje/AkeJUt2yVhtEOMufBc9LtnWbs3rx2ZPTwswAPi38f9JOula+AJYB8/m1g14Bk
bSp4Ptzjs9KywADnd0OLrQC3SqxomcPzPmgbH180cRhkQeEOjn321rJ/X3N73Xx3UqSY0aQ86Ez4
rJyQBBNe6h6PDygEAzey6ZyVmZ9p97OdxGA+lAh2NWTw36vbxec4hc9mcV/mtkmDyHZqoUfd7RHx
vCOFkFvn1GXfaQJ0wIuIfQtnqFbqf3YgZKvBlYM0S9CeEcWw4AsOC1F0IQshD8uwio7bPHd0Iq9l
HdybznBbeAKU+WlwCfRGo/OqINmYcqD96exW2WsyyXmCr7o8uuxeXd7OEEwL4QNAL0/R2YhkwkTd
O5jcsjKNMuhfx5N2uGsShQBEwEdO6QZvNLaCIgz29w/GwWsH6t8XehDGKRf1SsB26ADq7mKS/rFP
zUOng9kpNqer++2OCaN9zqO8Lt16EDYB+qKlA59etn2MZLD28PtxSTUTBYw/z8B+9Np5c7szvZPf
TrtVp2ZhWo8CpD4pGbb4r+3sDwYyti33q0fI/Rw5xzU/1gmRyCDRVQV9VfBl7yuTDXfHrJHtzVpr
8saQcQ+MSP8XmaYE+Im6Pz4pT/1QOOWMT5olSFbWrbTX+5tkr15Ot3F3fe8qrm4qdUK1aMeQTNa3
yRhH1ESGIxvTdI4Vyi9x84PnnqLyMoYs2zo+gst+Q3v49cEfzMBwMZ3T72DXdUVH4hjIzv6AV/fB
5d9DOrJVTYxiPxQNzSMHbDhsbNaQqSrYduiZbQ1YTs2dxEs6G864RFS6PYESMO8p3NGl8MkqINN9
BvPLyP27laHnRQAMAOVwB1ozFsSO6EYBIjXSwRZ0UZbZAtFmpYKvn+aOrSJa6D9DzC+YuekFbR/X
9mCiGgAP5nNtMzLF9K1GIma7H9cUH8fgY7BT4ZdCQUKOycxgb87ZhD0bwNSBj6mpm3IBl5HuETe5
omMP+bFYoAUEQghzf/hauz5BTcu8LS6NbY/16mMYRJ3yBA17V18tZsGXKO4MDVNfKqkw8RWzu7pP
52CvLJOYJNtW+DKyR8ULR+xQ9ZbGThf6xDFkMp93h9IU1WVvQ2kWRn9zJUBxUCR/Cvgn05m2lgup
iZZLcuuB4LgOJI71KBpV/1Ksmr5JQJ83FT2LmOkadZw+2VIqQyHwPVT6XAc0QzsDK6Sj6R2V7Kbk
EEd2JBibNJURWVX2GCeRvA0KpHEVrS4sy17hv75dfn0F7H4DlEMzaUPLL/nR+LWpNuhIPO6dezm5
MnRSR/Rs4ildQtvJIJUgw4U/WYu4N9ebqNsYm0o5TlWGUlvfwj9J6m5DbrO9Iub0VYMo5f3fBJQn
V+VVtxR8k3Y0tiVOOZSeeQd7BiUxioLe5Y8DIA6TD+3tyjxxwkYLgowHUjHkfC1YyHOyBhnPN7vk
6rH+K804d+5htjUV9xc3HGEPTinS5iau04q7p5T4Sf0GejO5bqlceMBQ0TZ8zbpB5/Yh5fvjWKCu
Tgy123Oo8kRbLe3pic95gX3bvGBDl80Qn45TChD3FWUPv48C+DLqGUL2oCW7nIk6/Ct/u8XrCxaX
urOWkG4D9pLnDYf0s9cXICXhhQUoCs+7TlWqHCd1kAHIUws+Mv3JmspS6kMZ6wYZilziF3iyZG6O
xqIFZLZqO6YrO9I5AD08O3IGvhym+mBW22AGcBaw7IhYdkv8NagjqeMvc5uknCIvaWywsptiW+SN
oEacOkYnQgCr6m5yaKDufPMo3f4X7kmVcO8i4cRNDoFVH95sTajIQqy3/HJL2tX4g4iRqvG1q2Yd
U6kbwEkzAeCj4rJA/JfLIW0eA2WkOzoXVFd/Cxd57NUGXJSjxtsjkCXOcmFMjF18FpTEAY82wTWE
K6a4JYcB0TpFejDu6y/OPvqE9C64bTWObsFsF5wZs9neJRtNcChrVbOAMAwdBhGpqDLGMcgcfl7Z
6lYK0khTx0dNpz7XOdj5EhHAeVh61xtz+0eDrAn1aFgNlze3haQWVtO5UHuQz1j5s6y+w0cpPU8p
qNlaYQ3T7bfISRPpuuJX5Rpm/WBI+Y3ThuWPIEa8wkRjB02ztXvUHwg69KO74r8e4CIDDsC/sURu
GjZsuhg5xAdoKSiqa4RdrXeetpxmN/Da1LEJjKlPOLHX1A5ViCwddfsvf80C/Md/BhfMqdMuuX4m
0GB5L1dw1y8HIlYMYbPsu9MSTOzcz/4+SfWTHBFnutccHtS0Fc5+dLcwZdmjdJSszZNqpZOgWVic
DXxt34VNGTnf7nBE8DmF2+Fp3OdXteRa/VIulJNsQ42CXxTIjQzTPs8dzjKXACfITrYlUrMNOcLX
xg/Gw97PZv04Noru/hsJVMS5f1rQYJ7o78g4jfXpMrH039K/X7FPJywnCTQsRHQPa9QVvtoHX69v
zidcNqpvK4U5Z+wQZ6LNHU75UIKcUXc18n1WO9oK8lgsD+hA2rVXBQEEER1pCQSt8JSOLK8Ik3sY
TW5ZwNFBf+SfLRutF0Xw69Zwg2N1FPocmKZIgWkG8A9XX8IJ0K/m0RT2oE8DvhsimVZ80heZKdHm
hn06wbJNVGwxBzaSI28tf34Q3Mw/UJOPea9mz16/jjwn5oWRGmLf+wEpaUpuOOBjBmcbvho5bUpE
BxCvfekxG6RQSWTptprIMnrQx6T7MOlyfxzUix+PJjnu0D5ykpQTD5QQXz5BiOAuV6DNUotC5zgr
NQc+XzUNXdCW2OftkFvtPTeyViN8GVhOHJdapmcBrF3HORmZyBq1CRJZxJNG7nLJwgiaYA/9yZ7Y
ftPiv/AZam3AywCpeCG7t74g7MuO0WbwuHPOFgdsTtaC1lHJkWN9hX2rn+ZkI0dJCpsN8xWJBDed
KEDBGt0iAaCNAVBcYziKzlqshcVsUywFqlMPSFdsq4PpcgiL1C08TLEDlcLBWNXgGIBY1CqrglHM
M/hXwyBL3dG7OkH3njofRpQBGBmknGTljJTGl4P+5f690KftF5Q+Uv6Ix/KAC6dIS4Wlkxo1MR0t
b8D1A3zSgS2OQwmozRk9TMcBKh9aPs90c0mPNjV08eBGwMTGl/5CnjABdCMKeLkhZcyckNyeFOg2
ge9CXaMwsp16FkPJrlKxr6zsdbYWaO3yMxbIrk8LbiCP6RwC1E+IGw9ymGvpvDRiLzIfbbOky7Y7
mbidC68aKwhgaJ1Ncc2gIG7t3UkbHIpeNK2ktKwAyuNVGW0wTOhcPML7SDBN9WRbTCimf2xxpgds
ZYSQ1l5nAaz9Rxdc3rUcItV0BVwQf4m8uXgaNXkb2x+2EQA1aOyc2yboGbZFreUJa2VA4npEnz5e
D1VjCrYQ9eZWOjLQXhaOeROY+m+NXhi5YwEZCDB1JjOFtbn4xuPeb89c+fNknZhD9AW4JVpn441g
k+wDyv1v96Rfs9k+6UXxivgfbahUG4f2WJ+4nAZkbC8gqG8knDr3i0D+hjvatV9eSY9LBdSawhuV
+aDxj45lUzvW3FiJoezfn0RIJb4NL5dd6cz6f8jleM4LFnB8cfYcd+y3l2sX7uw8DBxUvsFQxBXk
4wAWDZHOAyQROAqhw+LaMhEexkdXHExfwvGy5bg61BNA2pZA0AjfjfoG7djAxslfz9CaNANEQyNs
0F0VHaoGKAEam9Yt1QrFfodGflh0317ofiomsgqm4sFPP5WMseeLM5LCrSypbBSr1TyLgcvB30c1
lnpcCRZ51g/ZP0ItTnMKc66L9Ed/c5N/Nqo3zYfVASQBDeweqZnBw2zjHadtkEZcWT7Xq10He0NH
omgbdzLriA4unX08lNfUg+O5QwG4iJecsyUYUJv/+j6T0itm4CY4QGF6IBvNSd5grQ47gLab4PW0
6OMq/7SvWIbklB6A5XFHAubSHfi3JcBQhcDJQblwbvHgzLksxeJts0OzykjQ20FGgRaWYEU+GUEa
XKIqax+y93W+sTZ3pXkBqDC97eaTERbNUTslsuqDjqXbgryBqt+3EfQD/27ETmeB5+AZ57VUaOus
3NteT3IXw9YYNFYgdtyj1FJc2lz5s4d9cLQyg3p9qxZjdZRECCvTrxh91bkJotNdfQl4zL+hK9jf
ry7Tv9TaDMUCGioLwcnhs1qX02xW1ccyhOk7Yhku06Hnz1SLD1AeaaVd1D0UGwn+a7WclI5WmIJQ
2bjhwCzR/ai+b5nQJkRo+jIzhGMCGATU54KILDfHVD/hPNIIsNTUWjMMcQsMCoARW8n/8g54pSMW
RtphDTj2ZBo4mHL+f/GhVfn9EpatgF2/ytYzuaK957KP0y8sNb+Fi712iyv3f4znKAgOARcseqU/
HOgREgj+6SJww8Mt8jQylrsfL4e+axfvr6+jsA+445Lavd1MD9/57vagfPpXZhujK1is3G5INmBq
ZbLB8DVqMb9dtKF0zMw4MQw39k2/l5oWwZLlTQdg2tR68fGOI8p+799AO8r6fQXF93RHcFcisW0t
1TyXBSiUUk/CNT//3KHmT3txEcZd4g5cIW+VMqFMKRLtZD1otqRfw0X0Sxgylc/P9gFZh6+4t7gc
DAEm4HZdI2fYLJUkBsEm87c2Ol7ICuaZVkKdfFqY7XbRXCNVZQWbbM+SM1gp9xML+C7HV3qLbaAb
pxY6V5jbnBaNtWZWGW2BnafEHQrRFXEn390RC4SKYFqh5uddrNA4Fv4QGSWZX0vsiMjNQXrR6kag
nQYXyUvAj0BFmwMcUjDhT+7msqR92X4EkCyXULnVNtRCfB0WL3K4GB7I+fQ4H63tpHZ/tp2Cpu6f
hiqIlkoCoLeT3jEF0iA3ZyhQYlg9l70BgUIZleM92lAdLqbxfj1TIqT6EvTOrHMUtZAz1mSXhYcC
8vC1e1f5eWWrMrk/TQ3v6MN57ZUfPByfcn2p3vKjmhacu7WNQ/3xnDDapd26PC9x1v7YAokbosKl
FuULMHcIBS68GccDGxDmgp1cY6BthjeZ1IGjcl/EnNzQC7w575nYhRTvq76072DkhbLDs8B1Cu9M
l3EkcSkgpyGHn0pQBlLh1Y9XsV+YDESY/AVrCWSVxEAQupAwLiyPCDafIpRwWIIj3ff+hrSaQZsZ
0rAOubsjehyAePPdwK2uR+fJX59JdSbOmp13Uwq0Z/U948e6Mj+A1hUV26JKmk/p1yuqVKusU1Gv
GttjnzIvhyuI1me7v+Npf+V1tAT4+TY6Na3AqNhHMMQGeKHuBWu09JPY9FD2suc+KfQe/UDoBz5B
5gjGhZT3stUSAuG9nwwdjjfcAaYO7iZiUOPh/uCEZJ0502TcVtO9TdK4uyuPt1jyZ9DFezemttjT
xshMb6IhCD8wySU7eqgcop3CL08oR8eXTQV5xviez6t8XbltaDB+clpCRuTtQTDLx/Gs0bxg6F5I
DGL3Abk8HYiNMVKFHQ9qWL7jsWNGXADX+vmnZ2AdljzcJJbpeIrY4/oHT11WAjEOJT/ykKqxwBIx
azMzQz1FI8ug905r/aNpTTojfNdWbgIT0gu8LYQiZgpynBqgIqcdA8GLQ/DZoLtdUbwhaWBWy8yz
AQh1x1jlgiT+0mFoPJA1XoGS3LnKsS7JNIzWGhMtZycar9m2SMbfFrFtGEDcP/aGWaguBmQlCxRw
lObdmzAG15pmVxPePMVgQ0NCC1faMa3JU6hZuxuoK7WZvCyaL3lEhF6Ysx0Huy04vdjzEYlHm9jm
PFK7kDGOZRM74o4e7nIu7uv9r9uOEWPTqcMJ6mMhyXpRHMIsL/flxhQUyCd9gonKvNUgM+7XnLiW
5yFT6xVeOQ8jdcsK0zl41oHz50TG9YgK1EYU7lR5Xuk0+BxXcrOo4TfzxnPqAEtXnMy1SNRlHswZ
ZhCeP7onI8sQq/Ystdlp/Ph86nY1k0QbniAP7yHzM+9vUSm7FfiGEt98pxigKsZ2NQm8zZntGTew
2C0x1k02/LiZG6Q5HxGh2PcmwLi+eSgQSEqnc53H1DX0P7hjclLaawmw/E5FppxQ+NhJj78N+TOl
NmcQ0s72AY/BepNo5/+J50syPryT8ypqiApdmHcuOe0sP6pFHVPp5NSJ6t93ns9pkM1Y1QAYcIfs
pI8BBN3csuqkbOCPjDueB88b2GmUeP/Z+TpXoIyyeM5xi84YJNY8pIvjIJh5kgOFkg+E0psB3Nwl
wfps7zrrThDz46m7L+ncXdg4OyjTb6zQlefPuGca4EtCrXwvQ9vdqRkGrSvgZf+pGDZ09mM9/3Wp
A+DFAoQmNi0xQpRrXGSb9xkHxZhMfNu8RJe3V+GDWjt9Kjw7l+mq3yJJODYnlHrnHjJ0eBO8iuKK
GTtnnhSQJC7FgHAD3YD/DZjYpmr/OJt34VcmILcVK9HuCD425O3tPnslkrxQkP+xvRnS2Pm0PyYe
rX0+fdp99bSdgxO034/6AIs5sLbDWbViGaPEG5rJUUespR0UNTczBqlzjYK/OFAtTCVUOPgaw3H4
33fu3wuzr8Izl9B/oeKWEJuuYp5bTTATwRt0TUnQtI6TdQm50j2sWpGdKnZEBqelonhcJpWAn3rF
/jWhKNOVXm+sYJAnGlr4KGS+b2l+tqdqXCUKO0W+A2JpUB654htCa/NDBzXRaBHwYgUXVRYQSGhI
K4LgFvME0EekPxHVR/CgYsqRUeST/xL5Sob0CbDWypnaRrZqToR/4bb4X4KBIC3KBZbn+USq/gUo
rfY9c/LSaX1NMmyxD1shxG6qZz6kGG/NfVV0MgDJoGfb8S1za3CFHaE82KgVnJ6S0GZVivLzSp3S
IcW+kImP+8afuYmBR7Egf67HlIsRChtSJEdsdtTrkAhtvf68ynwRnhOlWWatr3nrSifNstngS4Fg
+7c+Fu9KRPgwjr7zBlV2UGmUGw77nEwFjdbPkovTrKurfa+oq42nUPVAuuAfSbu4VdGeeD2YDCJ6
9xATm8+f2WF0XSZlR2vXMpmGEGE0+Pe6i92Asy+xc5VCr621K+QAJ2QS2pa2zfYC+Ufcu2bUOVY9
miiyluSUMGu9Hyr8QDH552Eum3EvfOuvXeB0vF/rU3yMQij0FG+2CBQyPLgntXtUyMwP0f5uQreA
MbTUcO3eneu6JZnj5+l4guJYYWgoBUsgyrqwzAZuknZ2U/SEYdKtQ6Q0yzROnyNd6H1rayQNIDQx
btkjkTlQ3/a5AIegmluqaExdGHl550iB1kqc4l33IPwvTcBh5iARM7Ykoly1ZGTHycLQ6qm0jas/
skqoO1lCIZAa5PbUZR1c4Pp8k3l9UWclwwFyKAytcHUKoXGE7wyVUf+MhTqcxsZC88H5eR7aYQxO
6On1XZmtna1gnL0Gm/GAHVKZG1VdltRvKX0FwVkp0pijPPJwFWNeFYWjtcpzegSeyJ/NZMJ0XrVi
Fo+oOPy5SrkCVyktvofsg3rHJM1DkSqsNIm9sMWBq59t/zCSD3h7i72WUqa6IZDXdGmURYFw2iIA
/cyWh1OO9OhXftzgpudP1u8aZBIV7cbh+ZIDt3h4DNnGaYFu1iwWLAVJpBGKSAvJy0ZG7DEranEx
2v6AL8X87piIzzS+GcxrltUKk/2IveZcNDiJRpGdIdOTaO6V4AhXN4cb3MBQeVQAniX/rT78X6fD
v8dktcVmCrIVvJ6Sz73othdAZT7w0X0N/estsb7t5izqQ+9tqhLMmYWG+7nmCEaG1cbZODdhR1Cx
RPuU6Lm7p7UjC6lzp1heG7tDfhW3kXk9l50qYAvjyR2LnhUvfcCBel591bGJvK3Mdfqu1UZnSEBa
v6W6H0nWqR500V/s8DXkTmCICsUzlF9LnjOTvt9fpzWOcWc7eCxfd6ZnYO8BKObwmCgXI85vj3UW
6NkeCWeNrO859q6kbrpuLI9RLJ+jJIiilkbL8bD0sWokIP+GmSvPFeFj1V4/PyVbqr9giotFTte3
+tR8tOgD4sAk02dm8ZSCEjBC0OGC3G58z2uS8wUW52UL6Drydxfv1kyxgXElHRb4EZwObHZNhPAZ
hRhS1KxtlHRCjQmlGqdxdnJJytyxbPMFlSF6s1nV4QyvDh41BIOUcfKddmSxAQcC5fZevZ/SBtz4
Asikw41ur3odFK0U5bJKFBV0KoCsZhzZTsM4FlMhGDIxTypWu49gx3LCe0BA7pTNnNIDPYPLg1oW
PMyOIT/flDztrRmcw5d4mV5s8CzsVaSWlIL3Rv/UoSIqUYQaGnNSs8Dmpllo/bq5ZUDDNaLnGGQM
VHgozEdozakIY3BvGiezf/UVv86IAsDagqsFz7INwM9Kqe5OYdiesmT3vNOg1mmFDoCKDXRmjECK
NfF8O1yvcwUbaFHBLnJkJHrCMz09d//GSnR5rbTwbhzrCK6VlxiQKpJUfg9bC9+Lk42OMb/QsocB
t74Abz/agglv+olWsI0+lsbXREdN/tMgUBfAZwjuoVMbYUd1Q41elqRI9V64R6qxBthkwfcAI8xW
qRRrPV7P40JunfIn8RYRelJtu/SR0Dk6nXxvXevKBRdcaHklg7XLvKCeC6UJeiLsfB9IMih9ksED
/ABp/ud8CtFkKhwy3V2vhFe4JyDTlxo+ssDOklH1LK2b5bDQF6PV4bV707csdOLGcQSmpMmT/YYs
BO5uPR8Ku8iDESQJoqC9p/OOsWqjlRD9hi5SPr/Hd7XbN9MrXgM/iUqGXi+igXW1yn/Qu6dkvPub
0qu7kR6YTzLCYj+rjwl9c/CXA1EPYNPHsjZbYELmEpwQPdUbXVwrXWTUPlowakJxOopWjm2yTAAk
5PHMWJEstVp8uDuhLanaWWNjR/8vDzSEd2KFhMzmB00UW/wVLsYj4ZMB5s8VgqGRaeUKdBdso3BE
QQWO/xLJOmGU7wJkPsseKVoopt6C48TOCMJktNhdktwqCs7RftjI6UPRciMRnFkIO6Yi/ox5abmt
w0vITtAPHDNZ2jVmer7l3lpigOwYfr6MnKRbU7vW7eSvwiRwCvVw3baxHCGxioTtmXEU9k3QiC8p
OJVXSnq5fcXMIrdd9I1Nqp7q5wgPhuG7TM4hxqnIOsUyuw9eRuc6bCPH3GAMsWiKUWhdwLg9mCs8
G6AA0Qz2vb57cMqJ8uk9bpQ1PgCaOWNPNd6gXxG1hD3MsdE0VSbnaGO7SsJ/N9oIsJEQgPKbPuVq
hVroiZhyYUI0R0MppI9Osmj7h1eCbGN4CS7CnNtlcosky74GdTWsxLCJgJZOt7KcXTnoMXxxhLF8
G+wKqWIt31pb8I4D8z58hwvewpIrnq+5Mz131+1RGLFNPJiYVbGb73arCTt/pB90RoTshSUq2z0I
410taCCYw1mOEXi6IgmDWIINhJPIPWomRD9UqMLtCHyj96RqnP5hW/QvGo0bDO+KTTPyMsa5e1WG
lkHQy1PsnnmmPUpf3Xjk174KiE9dgZxm77hhLzOgl7PbZ/mrR+KTfQWgmBp/RJ5FlJA3E22UR9zv
Fi8N50sHA5GLI4dCMj9rRC3yzgYF4fygnaAyS2M4lYjYxEXGjOF1cjFBUfjKXGJY9Q3giALSGNlQ
YYJDBPlBnve/W4OiLEOdYTGikioRt/YvMCQOA6+ID+oH6C/i8Mj3rb0dpYphheDya4O6Qt27Pt38
wMwPdRcUkhlnzVw3n3Pf4ll/fdEiH67c2csqhIyU96mztux0FRRFo1rBGnNtx0H5eqwn2PtIWw78
JPCD/Jrx/dODOigWRptAz5O78RL/75C90Oa2rPCX5jNCSGkg5EVKkTfyLNqasvqi5OO7EpyP6GXG
vR1t/j9Oxq/74MricLgs8FuvIWdHGG+GE6EpE/BS9zt332PCNB9FAC75jaKajUuvLXq5h7BN5fOJ
E53JU1SCPiyezitl9Rm4kCmLdTZaWVSkeLGLcu9ht48rzShMiyaX1cjKhrMXpxhykMdMDVMbfFVv
vK7p8bD3+DHP98VmDfW8wguk3cO7WFN9yocdy+/UBgyPp1+/0v9A2KvgN3s7BEj9IqUzbFFEI5QZ
dEcjTo9vazDKq/F9HRk2DP6a4/7wg+3BAbM0AT46IIAgw+9txqz008VvgCbAkWOMcyB3r41VDvh2
siwTr2vPpR52ze24ET9qjRsKDGbn7omX7xR0l/q4qv5Q2vuuVZThCj5R+p73FRHi1YGm+G7X145K
zfeb6Q3t6BdcAas5tLHO2aZEaJHMNF0rNult8hGYxHo0k8P8xewva7o7UTTEvQldEvb8n40vI+pf
Y86aYN6uPw9zTNZPmB4mqZ1+ECGzhrZQurbQaTh0zheVEpVIawOEyvn3z+sIQgkr/vC5SGZuWT2V
mDWjOlps7qNt6LO0VdXac3WvdryPj/C+1IKWHaEzK+82vzQ5jIT07rqF5iF+sYaPKiOIk2rPtb6U
K9wcgVFj0hoqQdAN+/HpZsdwjcR72OHNhWpku6r1JGs7W48muuBCJUE6tyLQeLfVOayv/7gIlC1V
GNzSS4IDymYZjQn5IbCqEUIMVtGlYcCia70VsCat10NPPxUu7EZyiHdyTZPO7wwLL7aesW1+ACrZ
X0WMnepI+ngxnE5Fto6nRYYVsdLj2D76+wwfAbAoYxVxCH13q3bdhTaAz/L9TkrTyjnj2g4xSWEt
mjahC7OHYLDGNJ/9olbZ+FOfi4mN6CEfJPdNlenKiB6hShXbgHugkObZZFnBirZmEd4KSoMm9WGd
+eLSXbCc7cJImqyfHkBp79be2z6tlucbXrnwgQdHVE5AbqKVcl37wJcHccCQPT9U9CcPdsimx9HG
0A5535lW6s3lceHf1nIaS/FEcD4bbYPFY5rBnHJCFZaP+/zl/HsjaKT2/WqUMc+yLug9ZfxAFU4U
pYL8/mbLk82OTP/PRsvRVHkQZFrpS/iNFMwijNIn1PSNjz1Z0R/l5ePhZrG8Eoc2+cYXd7Qvm2bc
kPelbr85gRL2dZEasekDKsybDOKbPtn8Bbp968PFMfov5MKCn7IuHfgyPFPeLK+a5sxe9Dtvx/7a
rg715RO4eEBnwW7X/dMy82OIXHxRR4Gy5P7ycB/nyLm5QfQGKw4b7t5QLm7mT0UFe26kUNk8c/A3
dQPiQkj5+BKzQyzAyXLCDiFquMubMVx5yBHqxOY6TqAfiKDbINDZv79GcS7TL7zQjc1/kGSxPKyJ
XJRTK5sseL+yBgaFBJOt7wi8dwmlkq3LxbVT/xOAz8PCcX5dx7IQAz0rpqxtjb09G+LRLPTPNG55
cfGu4H7cyLTKLCFvfZJwq77P2YnVKeb8LRjCO9z0vKczsjdUsjxSyOPUXoaBReCLpsdzu6XCEeTS
UwB4w7KPaUiJk4tssPmqJByg0QC8sBZcCI2bl80k1AZc0uqzYCdQYvUF6VLy4y+6C42xn2gPZyXv
BHgKYRGcfSq62q5G/JFS3ZnOFo+INRZUXSgsIy+sC1k/YFfbU6BLGy+1o2q4F0y7cI9OXPeXCrsx
EUL7BFXxvcRHshY5z5N/I+k8n/qXvD6fCF9AotYbdJEkfPHCjuomk3pm4+YcuGlhT0ShucQ6bQuI
ljh+RkEE0EZJPyyoajvwRNJ1mgZDEN8fdO0yUM7qnQnUzo0/9nx4Pg5luJsSO8nnOEo6TDxgborh
FQj6nStCv6NAMlJb8YjuLH8iw1eFR3dDM2VLahBsgTdL9ylLrBJ/n68nsO69FDKLyWmtjkdq82XJ
+UF59MEHzx8k6+IhTiZNTDwBY2rVmwJFIL9n6pfyWY+5Ou6drmNf/hsnViOUNLZOFqw3YvENU6wP
LqvosWrr5VnizmuzRtMIrEvNPREMJoEDcDawOuMcQbBpUI8xFddJ+7I2PzE5Opl2nL3smq24IvtX
Gx5/S4eXgePERDScSoUt2WM9k8hghQoRrQy9Ayfly9HuMdLA5ccAjw20CS7eYzLheicH1jc4C6Cy
xoVXo/RQDFbzkkFqves3pxzsIRSj2vZs2C2Q43gEbtzDndOWevWPSKdNd7ZQ3bDg3mYcmyj3zjFb
awsc3LYqsr29en3lOkQTgTfKvNv21bbZW0DB2y7Ks9EG1mJsuZ6fXYZQYA8CfMXqLZG5J6ZRmQJf
+iP7Sg4iok8O7NkXLuo59445pi+Q9Ci23lMgOlIOp5vCzwAmObZeMCDa8mRuolr1mWRyGAtV+SDf
XufOQAN5MvBEcq9s+W8ss2GgJ5dwiPctNn4x1yjdVBqzNCXdZ0fWDL89JeUnpiIxt22mkEjZWDDz
HJhEntA+MdGI4Roc1ZchR1v7eSqLQUf3/TcTM6Uz0z2nTZ/LG0sowgEA54X3fWDiWtkpnCP0odgw
FvJeXvAPQBCkMolwWYYLQ2p+BuGepS9kkHZxOlQSrWaK8xXAOYwxPPOg5ipjIIBx0J9feApp8Ai9
vhwAJtGacLHtxFJnEtnCZk5WYyp2TQ4G/owwIMhOzmjmWxXqoSRfJ+hTXLkYmnLwiIzOEcPY+Lv7
J89kvNP2iwpLhqwyMovG+Z6XcHMbcQyOor0ZnwEwvkK99kU+7oTBTWA6OWCpZYtVe2DIFPmoLuBr
iJhwW0FvJ2wmByer4+lJoYizSh0nqBOy+p9lE64TKbwCYPgkQn9cA8BaqsWGbzZmTFq8uE+E2R9V
cT8P2ivKqUyMJDKK97XNZu+1gxH+g9LqToMbQw5P5fXX/HKwOuym/pqHmEXyADOpEJQOoEzJ4hwJ
qVhzakVinLQuJ6EXVN4VKU1HaUawK/0jdVTPQOwpQ1Gs6tMAHA/9mYEtkRnrSi1C9M6w+BFiDhdR
Z5Y6sTVPa5gTx4KEb2Evo5Oy57UYHEC1xUIvek/xYHJ2Uec+ph/eK8kIz9aFpE9DXTwZeP9g6diL
fmtgdY+imdKwwTEzRiomZKMWHaCnFOKuwfoerzLVECWtGZXxCUpco5iqQEghVrtBK8lg9nPwvNFK
gnm0Y5hkJBxUzoPNk9oA8E/7PlOLYVfgBAyzWOJxfitvckkMMq9GTWY01sO9CHWfd+nLUESOz26v
C4hzIU1JcaW9t0sXK0qbRpuwhsc7xYzp2JtJyxTU5o/55vie2kLy41hwt+dcSdQIE3b/JFdCal18
f210tajc4O5xciasYR+2YkOd5qVyT/n+0bZ7ZrnLWd3+1N6d24F8N2BdhxDdCyrG1wT30oqtoGAS
MwHK3j527mPCENtuTgDQhC/9/Pb5dC1kOXGFYrQngIl9ANr1G/8Vkd1vXBlFf+amYcvxiZi6KvmO
mW6W7C44TPjlUSlC6iLiOxLE+xtMI48OYv1tHPBeKWt27KrTFVAdzrSuNwvIosr9DRJAHTtv7zim
/gKNAhSaIZThsllk9dHNJSrYCr+PTNKM/xBhElHqIBFS0dpX46REhqq164wCCD/mxrHyKZ0+P2Ce
ZwMcUl+kbBUaOM0nM8BZ5Ky4olM8KshS0cMf2kTEf53EZY2u5zkcNWL0C59paa3fEK9BOf8RtSfb
Qe2rEfPQ7lMD/tfyeSHFv4JxwGLUU9wqhtgp3aMr/Hc6BtwXbx1z+V2vB97ZS2V5WpWLpMDRI1r+
V+9UplAG2V9JeDWcz3baijSvF2rZDe3jG+w4hWHQmZNW2J/jSiGf67TPrRrJtcC4d8gvlZ+/ID7U
PaZSiD5x5w/U+d/lE9pYrDYTlpIYOmMT+Yv9Ou269WWRf/6MAIChELjJycDQO2OOm5nju3c156ff
pGr99i/qfdf1LeVsMDPn+K5q969ImFa80c41gkGb3bjKccZ8UBw5XgzTRVASJYrgiNqnnAYGd4a2
oHewxmpgukT6ex+qzuXHvN8pVGRK2zlX2W46mGIvpqrX2VWSIGtVfccFB7W7HI7xoDZKai8rBpXp
5PwPWHb8F4CdNjmkqglhHnv7MdEb4VD0iy0rIctx/DJGY5V3nEKHDRtLhAWghrtB7XUW8t6bfmhD
rFhlHdnERu1aWC3SjuFdwa7BgD5bqpmEKER0lEhVagWCPZlERRLNEStbu6FZ4O+IgelVeggamwZ/
GivZYv1GnvJ2WYObyafhTKaaXkvtyvjsToUVCCvKmYQ6dwpqQneSDRNqFexPB6yzw1aASRZqUKfy
7wqxcM5BDknOIZ2oWNTy7s9ghjRua+WewXPHDom8PwFFoW1kapxtit84vj+LUDil5JUYRVDXkDSz
huHCf3AQsq/RKVsahgTa1QOzhrhJI/kK6j0D2iiGEl0g4NoMVRxlTjRMqY/EKW4B2H9sH15L9LOg
4RJxBu0VPUjLq/0idk73a8HyriolxiJTLu3fFI22PuAFqnMvxe1Fa111y2wXQWPW5hoNcV48ZUmI
+3LbRqHgL6O/b5zr/tvycMdoIBinDbhQo0pYyT5sFd+sXfcgT7yq8NcIcvLOQdcrSnAuPXSdZTX/
+ZiFnxlOrYdPxRciMRdKJZm9DB2/gSLawXqOosZumulrLcDXPv0lz/RHRrewh6wvm0RAGXN5vKtX
UshhoqdcCT1OcUsUQ6Ai+GgFJ6QK2dnKTGKRSkxCVFmYsIbrSImP9dIh2pURkxldhMLg7cbeB5s7
jJv6Mw1GTHNy+x8Mrf2s4uQ079OfFNN+G+1uwkR4ZP+u0LjDDnHdCZG+9DN9LfU/s7b+lPtLpyEl
TaS1pAUnDegV/DKMaad2J08XZ0xt/l1nDFbUUrejrJesLoAll6WULMWZGmYepJy+0xjey6Df6h/C
VsHq9TztayNU9zWIn/a8LD7mQhalFNA0uIMZAdOAS03y72VgeW9C/Ay1sj+IkuzRzYoqHSJ7fUZx
A3ZQ+71+5DfruHsEyVbggJOXZ2HX7Kso823PJFlqIB2Zpt51rG1UgmqNuwzClU+TVRzmKlRngWa4
7dXM2p1lVA9l/phi4T4woGKAqGkBmTzV+lMJOJ/jqvFXnaegwHMUIZVcn3/L8iJfAxLvSeM7hY24
LXqZwYl11bTwDNPzp/VXTT7HHXvmKZCQMR0L6KQgIm6CSjQ6KbxU8idvnmWmFH9kqqdQpZn7pY9v
UYMPd4fDstre385hW8soiN6nfUvycRc788QgMbCdR04eDSP3hn0DiXBk2WCPQsyMQqyRX9Dogg/d
DJtVsTR3hM/D26/Y9lgH372npyuhOvUxgZWGSw3b46B1ID77eHkzOjZKWlInlVbdTE7FN2BCLgrL
CvliybkSKWESaWoyZ6Pyx551E4kmnJMbGQNWx+9pYz5TCCEZ50bagD4S2UagXAv9cQhsxJv5RG6J
hDsThJRlqRJSbiQYYnfJLkXEsUTbdyxFG1623mK3gjNQz0hEY49U1aPRYVpSQ+PM6kHabphdtyub
lNotDFUjPjykwXThwQcSAbZs9gp7XyuUCTqt5z/3WjuVBPrYzfZSLQ1Ilzr813j4qXEg2jVQCsdb
ConTrQ5yVEnFoXEtZJTB8k3CuL70P7cc7SNRUYvkoZIGAbggb26QxrmZApX1gWaHFhv3Gjy42HXH
VtuKxh4hyZOxR6jDqJJCV1vZqITRSe0eyIPsGA1Wz0ivWJ30xJFwKGTXNpAFEJJuU4BhVEKUoQeL
K2NoeOV3aic7vWOrFYLInYve0WGtg7k4543qFwLh50bkoyDwGscxARAZulTVwfn7YhViQHagAG2G
5cyEr865O3PXdPBrNx6jQAB0ghV7u3SV5v06vSZPa3s+DW+NU4bKZlGugImTibItbP6uub41uYG+
sOM/A7alpTmruPmjcKAxZBqBsZUJhO9IHm8Mej+oEdvJKpOhjUQPHORisKqoEQJbtkkQ82vEi0u4
dCkBY32dWK1CWoqxXmmXnX1EAGOPR84+AjUI02pcQVzk+eb4xkuSNcIW+Vysr7BMULGhAihOcN1n
jVAQQkqan6Vli3U1b1QgSrYhITbmvEyrZAxySSOb4sKhaVES0+Z1jILXueeUYLHxxEMm2g77N9Lq
cwjcOpjdtKzeAzBSLmjt5651t1wmqDmT47CVNjYfSZIMUQ+LnYiUwuJuXEFveQSCTlfGNbdK0gy6
3Vc7AuZ/T3j1M1OQ+b8LnA4GiNY7y5Lbhm8KaG0IXZs9AZVJaj/itwmwjjj36aC0ePtas/nIsOyb
VyH6TtOeXIVUnwbZK3VPSxZwxFqAmy0hXGDxJ8D2b3PAyH7FxOo/l/ya9sSFRhkjpB8FNmsFROAs
NjLfDoUUibPAVXMBs817C92p7Jb9aIKoFVVWhN0KRv/v1y+XFql10k2YjkZyn+qirwnz+4qMKPLz
piDCBx44TJzN2durqQ/vofvzXEn3kRP7DEEIQbXVZLIjTymB803Q1b/gJtXbyw2eB1/PGAtySOio
BMJYDBHYYJE877scQVvIFyWs+foHP7FM0KWnIlFhh4fsZ4zwPfFZSc8z2UrgqSbzBZNoHOsJ50A0
I++c4CcT03XBcZeEw/C7gRm+JfTBrgBhQU1DGefIY732uwGOA7f+FThVKfyWO4kpQxGE0UCKpRyK
ue7QXbR3eiqBSilydIHuyFOpJVhE0NKKxLG2ikbBHv3JzqotCjeSTZz+mvF0b8s+JMMtlNv+KRy5
cNMN1l8kv1bE+ZnrqNR1ndvRYBz+ctshidxwjVp9NtH2+tYTncoAPI+lR2DqPeWSXKBZCO9iiYnA
JqyNQD0euMX7MULwmdHcHUqsw5B9GRcWPgxRvx8vSeLuDqSESv2f23r7bo4Ouszi81NKwOWrLQ0C
+7bE+3U93j/NswWgDFK2s8Q0m5Tr9qzZtW+R1y7Up1xrZiQky9VBrZ5FExgI4nErNwoHMmz/REnQ
BBn+XBf/UNrdUb7vGyyc8Jvj1dnK2OzwhsCtrK8dx79cxtx8rAGA10IWW3RqJWRRRcgBOWj0xh2E
Ll/uad5F7uziVhXJWhGdixk4nuawjkc/Tdpuv90+l2t43sVsvQ9F8JthzewAwvOGpz24KiTLKg/5
B1H+cXOGkz5ClDjc0LsRzbKzRchIAPw0XMfDrWVE7cQzr5C44fvGI60J/dgVXcdS7P7R8CDIAnyC
pA7yWd+1Dp2yqw/B/O2/UghgFl7MDBbCDJsY0atiUwOegpiEjTbulo/KIS1qqP/I9uhyL/sWTejD
6i+em0sL0aWVwCkVKtlE5+l8Ziuq6AdLP+xc/BVCZLmhk6+S6uluRMnA3q5OJRAXRJDIw88pBbb6
gIeJVs87P69+ANiRfc31deIXSfe2u6eEibBFu1QfIvWfeB8KkxURGW4aLiQozwGXKvgGbbnfy/kw
ekdnrh7AM7SjeRgaqwJM/Sw1Vwcnn6YP+WNNDgP54CeWWzO56sUqabzEZG7c2oz6ufu+cxRnQd4F
XMIAv7huP2C1JY++Gc1cNVuZI6BVJdci3DD0qFYxLjFOg0Qc3h5FR7bAu3DhQLyHIpd4xqffZnTZ
0bTxRPTI9KA4l7qYNmjOFQe6nYMfAb9EeNjLG6Yi85ths77G2uAxN2njhREXWh6J79xlh2oxSSAM
1L+kjiXZSRhEyVZTo3yhHHNGmDLf9ORuWcKjREtJbFW82evm0HuNPhhDVSiF3rQxmOWtLkIdZihN
L4sTZUYC7loTXYbpGLExZsVIy3xErw6M3UBLpp7As0MpYBOWA68jvDRD1oXeuawerqfkMgudFCSx
AnuebVFL+V9a8x5/UaJVTLn1SmvjoQsawoVOCoD8A8ozI4BtmT5nfmfsNT9yDoFvX9BfTwNnLdRQ
g7pjDaQL8dAA00S4J9x02uyxIxTm9GHI7VP617SNIJUKd/Ha0rWMF2nMe5lgF3YiJjy3AWK5eXpt
xCPCnHAmpM20wUK5+DaJVeRVDhmMbMtadLWsptReHhP64+WxJdXL8aqo0NgibPwmBzzMKE24Walw
vvKaxjlpvOrAmmQNR5OLV+r5nBEWkUM8zcbvfP7IwfYybqPqrK9EH3nuHQkRHZsahRr5umPLCKqY
SZejdc/Z3gjcHVfBrjsBods8FM7dOCmPTENQ74Ptm7eKcdTuKK81qjqAYUXbGP4X8jGBN8csJioa
BcqCl7MJrE/vrHQ5K1RaWE3e6sfNYUiwc/o71m1+EXLyuFh5ywvOx1obDYT3wex5RLDeD6e8bmeW
AZYanZdJQkGNyBalgxmk0JetsfVkygPNbjAaTefeDQt8n35fIYcg5R1twqV5tPO2ya1BqUa2MpCx
2FO+Bf2rqfkY0jMgmKat5gmrPBBT/y70E4bdU4KAnC6E2u47T84zbjJgYRydN2iDf1x2NRR9mB9l
3GpxDSLkEa7NeZMvUpc3KkgoyAaB90BKre8lF5bpiand2ip0tCNaJez2gCa1iiyNWnbPJpv2evr5
9HfSFoKZeXjoNAEZS0w4m+cLABAXfTWVjDWdTmX5L7iZ+S72q9wGBYWFqoeCxOz6SVhtBX77iU2T
WH/x1AaRkN00gr1JuEtbd2ravePyD882R4rJqFNhQ+AKxT+TTghQQWAMDFpOc5h9SlkFPLQZvKud
I3ScvQy41CWfz+XkNE7xDPO25CcB2P4Nxyr4MYjh/UqJ6kKaQ3wS8IXubtILk5JfSQeRKn7bJUFI
aYtifzjImBDk2GlRaEkC/4riTL09b7WphAsriTkmscywDNsT+SHHKmn0V4Vvg5DTZrLFeK+kGf+s
cq24S0w5Q87mPW7iJfl2K8+VtLQvulZ6nPWXcPLZXGHwu8R910qCvY0XwgeyfHs4sxI8j78igVm2
7vgmEMViyOXikSvOMH6Lfr3FEh90Qr7lcT6VR5DrHT+fAGgAvVLYV2LEy55niMBTQGF9gBjOZdDo
y0fvsJxrFx5QVHSJQZr7JdWi7qnKyR4HoCQe+ZfqQd4jFdgzoG9IE64/Kn+iCrJ+j/vZdMYvJQxI
k3l7VxUE+/oOEsnZX+15AICxXz+IEGjInlSYUos0txdQEQnwjurigGBA5evj+O4FnJSi7GCFOf3v
WEBMO3BDMKrCvL1MPtn1AX/JpgRwj2xbJlNt4/JMEvwvBF0IQ8oHptl1IH139GlusYoG+tOgc7JR
0aayt/+PotDKocEkgGEakVILi68mG/ApjN+hpt+JpK2k8IUbc4zcZpghA6adMnXV/DYuuoX+r2eH
Yxg1MxjWdFEKTeg90lBDasGnar2lqeEQ4P8nNFEznehhyBvcIOB2n9kMM83huqu/alpCRomUWbFG
SFaxv8evH3NUB8C7/XE9YolOLHvf19SCNyBaKEZF0LpjSAPgZDBzSG6nAy+1WFbfaLEqZYJUAaat
4d5JS0yMFdYyLM8zuyT7DEPWqI6+hNIMnYsVaJxYuytZEiuDFb7twrjHemxXwXD9wdr9lK4GIQVZ
ux7yokyINObR5MGy/HS0YppWXLjOYdQRw2GTQUurMqr9lKpdz3RQyI4nUkpjCoqtQmnxpMOYbw6o
6cECkPEUPJW2ErWUttL1sLnTSKBzE3x0ap7EpWe5TwPERvS6LksSrChN9MBjHXW1fqqX6ji8JO6b
bv8dWY7rtig/p9gb757yI1aUmCyZyyTjDxObiu4lmO4pdvVksCucav5qO84prUMQmaFqkGscp2TI
UQTOwIAbCNr3eVGb4zGN1g4wiB+2djJUY71DljL8sCtfcb4qYNDs6Xc7Bce3BJ4VbuOODy8MRbhv
E1Bn+6hswk8zaFTxU4ztBoJvVaflGqTSQPWo7ulxCGtyC5q9kycwJ0ILIH9KC78diWfmytWm4OuE
ecPoHhVi3SHN6hPr1+flPSg2Bjct7chi1J7iZvXZMpDBfCkcNghnUlhdmiZp/uPFmPB38tkLjmNZ
w/jFfZZtZyiyBdxgzJ/xGYNQmWoIH6/w8r64oOTsrIySs5/4/c3Y+3eI1Q7SdIk+WhZp8INeomz8
1Esc3qyL8jzCeytIhUclAVZ8Zj86C9WgL/yw34B3kfMauomh2wSosINcmcw/JDOyRDnEDxOHFRKP
RHoDVNR4WsikmpR+SlTAJOIerfJ8OB9uNfUUneFLIEQnJaJQmh40KvU8mKKh0dUVaZWuckrpKujg
ek9RXA7rBA9/ZktqKfutYxMG/VwnGPsF8oN+3dqbohawKxSXG1VCoTLaKBQck/duPIMLbzCW3bl/
OS6esVoA+1bUfnkGyDmxRP7fBXeVGuV7E3LywmRL0i/CWRM4lcg7PWGysmcUbymOsd+xgbxnjCz0
6pTUYNV5S4euY7QK72gri5QIsBucGcNXgWQdEHiJ7ma31qNR7hmaYp9+6aBfGPmuTRsZsUj9tnFn
b/zWbEmwGf5Pbinux4f89hqOkQJRKTVSo0GaIdh8OVSq2YbbPEF2lIitRy1eiP0BepB7LdlL2hLg
9cL8Ym0LKSB0fUpo/VSmR01rv9fsGBSaXuhUKZaywEkZreHYSiQH0mJ7lnFoe114tLA93M2oKgQn
hD4UlfyVJSrIY/tES6EMrRzU1Sy4M89s9u3bV10etm4W8rv3X7n4AjmE6l5eWnzFD95+3exSvcJ+
aPcNb+Nhl1MMKuRG5Y8DBHkOn+84a79YWC5bdS06TUMNbRMyqCVAf1Vhi3d6FguNYfvGICJnTiql
AIKsYvGEfiHa2A1WC4Vh/8rolb4rCVqk84nK7ZDOz5mXudxBK8z43hgiNIgJCb8ylCGHtDYOw9IO
gzqoyWr2h+AEMhWGs56zxRKYERw778nhcPN9onSOGedq7PLL0CYc3xctTZway8opYAcTAk2sG7Ly
GTK4hdI6KCzLp5QQh1g+Wt6iT6Zd60uu4289ZSN2M/MNnivUI4XTULrwv15DjsfBOdUlvpMpCece
DUi7nxBJvOW/vS9A39ldvOZjk32pzZDKx6yxYCXvq1jD8Wq1oJ9NGCjGgC4skegb/McZMHCaSGV2
oYskCzUSPndH7ON6VxT6ZkqPW/Vo7b2uoh35uluJVlI5belqVN6mXY8iG03ykKUgkfrWmASY25Jx
kCSlEhmtnGD2JIsB8SWm4Bt+r+fBN0pPHFbKp86cbEb/3GeZN4cYNIBf0NdWHDlhffHdBKhg2ajm
/9IINb3eb2xUHtUmR8dErm/nS2gZCC1FyaXo2kcmvlOIamjTiX/MBshKhHwSc7SoE/GTtvrXvl8h
hTi1M46zaoby2x99FC2PemRW+B0VItAV9yWOwlIO8obHjWiXm6dYwNbpIX7+Ro+C1zCe9scdPDaE
xb4A8hRSPhPDBFkuL0oIs2+CpgLl99NPgGOOBTxyNAd1VyDDpTtz4Kl+V0ruYCPrD8JISMYvw2Tn
o5v2wq4RkoCw+jrSJ/Jl0X3VzHddLCohJQftL+W6FbmkSdUputvX/SGaZNkAwphvobWBmT8F8rQs
yguaaNQenlJbV9GC3zLgqQcPznXp+tmAWHx8dLU0HintLXkOkifpcJibL0gR+ZLfm4ihhBI9tEcB
C0qbUJmjV3AGWuQVM2rgND8cIRGH93AlDODdHVH9nrPcd7LV3yztZktWx2dDmTbCtj82sXHrIxYT
RsTQ11CaLCPY5eaUiuM5L40qP7EAzKgkF+0c6oWpdmTDemYVFptAMpf6GXuTael3dGfTe1J98g8o
X/anFx8SXuoCOe92T6CjkIcXbkkSOZotcos387VGDVI9v0PY92l01+oV03SJyQRxmDBrVlOH+kt5
94U2ZobY0jYCw2XjLUztnogKOTMpFUbX7k43nhCND5B0ajSk6dqxIvxBV6o+XzMK7TsMXj+hPSuB
rH6aq882jOcSv/wZSooC/29KdH2g424eBONs4VO2tXFb0nK5TvCPBOd0Dp+ds5BahqhGKNCfGqEu
pb48IJy5UslecN6EV+IPq4mELfxiVYE37XZDRPkYCpF6cAeMTccKLe0f5uTEJaHg5+IB1UYpvzUO
CZCMy/c+CNBZjapP4u3KKFRv3vGUuO9Aa0+whXdQ/hc7kJy2xRk2EnJddE8KdV6dNmvAMYTorReI
rFyTAS6lJZ1F4MCIayW7zORmX2nLYDCe2aFeuhV0nw/XMttMCVXkLWxT1RtnqmTAmfPXYY3kPPC8
yCNGWilagAYXL+3vMmocoYDQ42cD7ymDjovHwRYwEjc7d1ZFht/bqNApqBUa5xzaeeiztSHe39lH
lfw+HddO/D3A/bVI5zav08BsEc+8A4FhPlJ/22Xivxl6IcgsNVNy6qr/oSuvC+FuskxJM7wV89Go
Dv1GoHNNRW6s+P41Y7KEpaVLOmRRnQFsznpVnS6HLajOEmz/G38zNflR4cpw0QMbBf4Eky85WK6K
V5K+l4UYGfFcv1baBXZo89hjWc1wVkX1xdCcJSmQmM9Nj/XdXVA7JqC6dW31EqtB40fRgWXcyZ4H
LbDKBFDlBCNa8JRxwgT3uTu3LIElGJJOZLvDSdEckakQjacGvHBVSGmwyugjKo6PUfCrlKJS1cIL
0z7KVv4yHY8XphlfOvv/hYSOdzYzVH51nv9iTjQoa71JR1Bja/GYhycPRyQSFjNTPuw/3NitF2Ky
pY3gzEu1vgqqn4Je50+/oghkjso9PhI1eUt82FwLuTt6ToAev52S8Md5D7EbuC/Dw/YsTBzZtshU
nbV1Qj8JO1o5BzWrFl27eonqbEks9KYDZA25T5n3oITa1efeBxcChbNgJYPuHFAA34Vt1XS87qJw
LPHunRwApwZzHWop0P8F2dMLQeP2mZkWJ+qH+vX+6I869AhkyZk/v1EmW4LXaoS89J2+pX04Z3co
TWwP35T6kfrjP98Ch9mEQHa5VBiEQ/1L3OMvcUwnGkEmjPQWKXe+4QS/vP81TQ+MoBIfFpAHT6tv
JR7YJfsg7N1E408aUXn5ClaQc9nztxZ0HwmftRB4QEdPjsBcacqMKpzWQA0SjDk4q/U6TXgrkHCc
UAMwCrH2sfxY3M+BmH5SYk+mZiEJA/4pDbypHzVDqzwLJhvXGWnujXGLcroE6ektT16tF2x3jKsF
ClvMO94tvoYmUnOnXRWwdlyGDgjj5/qhbQ6VMVA4URfXgkX3SYPtg9tMx1sO9Vtg4iRzD5tWqeIN
V1r4M00O9KPRVmq0nQZPmU9o+vJwzMZPPeeDx6fa5nLhbVLe1KtPBtF05KSgOGZDbMvDWq0Gygfc
lV/UZWQ6XV8jUVchuMXpPrLqUGDFLmtsvuIsAZPbwUwhIhqA3/oqGd8xiIsi0/Kme6fT9rnTumZ5
UGxwimR0a6lhvq6zRSthvSO3P/8SvMw0gEb/Z0Riob1sO/AW2eU4HTPfcZHefvX3gAxFLS6InUT9
1zfaxBaqDH1BHc+BsSUYrB9lGU1jo+cZPz4EhszrFNr5Nozy4ryXFrkxtMc6RQaq7c+m1uMBE9I8
UIcj0PcbmKzhcdAPpKpg47yUmZOphlnnlZnJVFx9jSnT0O9vfENSXuST12q+pbf7K/kjhX8P7H84
JQDJ8r/WT7L6Q6ON7qHi24BWG8zJZNhIRPrmyb6J/KZ2L+QETbmd9Ktdz0WmLU2vdZXv5frFf4tA
/ZtpO0V5EGogzFpHw7hkz05V19sQET46OIwkt1vQ2Ao0QUEgg9cB9ZVNKgNXFsq8/dsJZ98CjynU
MR3aD0cirs10sGANcHILogNj35ePB6Yf4dKTq+1jYkRSwAml5EIdJ9uTQ+6lSRHZiOWQ6+hCPKK3
Bo8lj4Jb42J0mmofdGTHjZAdC7s5x4GIhEYwZkP3GjjpY6Rg1DED/QSHa2at8fv4iFYn8gXyy5OL
ghBoPcSW1M35dghHXex5Oexs1TK/Hbq4tAs5JGY/AqMHfmlDldDtyHsSDy72Qg6HwInedtoVEdv8
KRi7+xoWcsTJRnzRtJDNaXZPtvMnPOv59l2ty8I9C/wVz/W6KzWaXt+a1+7DINZZ0NjmxuCgBGIP
TcfqsoyuiJ671bJsNOg+9eXXnDLovZ/XS0HKKdsNEO0ORHdFlI0aU/zhkQD7csvW/6NTJWceswza
eLGiRgRLE0o+h7+ZkKI/yU26YRReQFGE6uBXbqQLbXp5H5SsnIgUWJaQnwBT4jkR7pdf1y9m5eb/
whCWvDJys1nAvOwtM5WjnvbPxdaCtfed1pTU5ckpcP0vM8IkBwJjC3CKD6hxBtJXGVWGWTXwWH1p
99WI+LTOtbcCyYxVHVKaD7zEwjrESRbfiTX5uGSICrUwUGvXO9KEFFV9FcE6h6bNm+U+vnxcUApO
Ji3/v7m/cWwRJ7cEziLR21fJZ4YbUGMlqaOTVDKqrv4naFrUn9rsyPKwMiekXNEsDynrZVHboA9B
/lU/IlDJmRJ6w9FknUhwbtfdRtW6jtRvqEydq8051ENDiPKF74ieStDTJFebP05qneMK3cgjBy60
ZJuJ4s/b660FMObmCwlMC9i7vxd18NwVYxzqrSHM43FtylcQV1z0l1MkELS4+kUxyeGqXBeM4cdS
yRjmmNR2YwX52M+OIEyPUBgGLfevxWY1u9M6fXNkfzfOmMhlmLJ1t2xeCE67U2vhXSQVsfcdDOOC
72lwJ6RE3JA9P3ynD6nvcgtPglLOmHntO0yyJpTAGD5KxfDmxrpNQvzVLHXZgtXrwCQX324tU2Wa
o4bCHTQKMDS1eFNralb6E5KfgMgnoUuID2AXYTU/9R76VK2r4myQ8ht14yRJOTxdEDk6wGCSnK1X
XJjSzR6HLQnWzk/Fq0OvylqXWEv7p7bS5l9/qLL0eW55U4a5B4UQjE+BbIXfxOAG33MF3a8fDeIj
Lirpe/S4wtotShDzUZABN9TBWgp1t7jDWLUGzqKBaXN5Y0B2Are4QsLOFrPltOiyWqhwCGHBI3BM
t4awrbYh1deyNziKfalxBZhEzIqmHtrlIYQutwOodC7EPJNiAA8AdAjCMN49OSPnd2M++44VJMP+
mhSkqBI42knKuEB3+MSMqPpIc+1YGFfa4ns+9ukOHg5Hueb028TVvoOs3xEjmLzohV5hszV+fmLw
YMTZ8VlkA/Zdwr9QuSUuTMS1xjutw4vr+xcwy9E5RxM3D2QVlW6AnyrASZYHBcqj007+T+GnfxQP
7gjwwV5vr18HRfh8LrEgR2H/Fq79nSXs9TmC42Ids3nUaSkPIa7QhfjMEUnbW15gMP4eNlCQ8aue
Q39u7TkZ59YDK6J+LdJdnclCpc105CXsXohdLCMeT1Hcns1Q5o7WRFXrFRQ5UM01xp84MaGTxyaH
3COijUreuIiQGTE1C7e3Dqon/13nczsu7UvoWp+lqHgXBv1/iMwqx1S3knykjZFMfy5Z0BIs50Q8
LE2FxNMhUtK09Lq3SNfopJUeHtSM2ki+Zi74mEBTSVk5uRmUdraNZL5957SSRoaDtBQfIc/r+vwN
wvlWqhQE/361duxZzwxv64prSJtvajuTaN4EEjs+gCqlGf289lyevJnJgBB7DvN6rlNtprtSd94a
ZV9uS0J69onVGEkSC/rL1w/9spAKtizZ9EzaPjZZAPKJHed+YtV5Aob7ti3mNez/BdQQZSZqjd66
bdrVqVT4Gal4UTbvg+fPwZzAzYt/GWEPgsG9sd0jspQFOrIVyldoRc4EPdMXwDmZJlT1gGn28hWZ
JV7Sf0rSSxf0y6Gxx9J2FL6UTK9IFb/nVBhJxIP9/43oqlSseD8ORq2FHJ34p68PGoHINhHSDnFq
mLiII/zGNFfg46IckW3zijKEqJ47UJI16pAbGL7H2EAn8V6LpazXdQGwWuwHmm1MDE7we/RnS/FY
KAn+gqu8qQEOWP52gwkTbs9QiH4kqqFjnNBbnhSkxIb0dNIhxBXB7MU2gaeVIV/5yA2fuTYCbCib
1u4f/yedUPg/5F1vTddUXz4aypIWY2kwINlTRYLtf7WrNUwC99BF+esKLfpXYzcNGZNvV5P4MoO+
P2QuF9uDqmxczw4d80E9d8WeOvaQxvyMWzYsIT+QtObxoGfRzXeIbtn5X61DJMbTPcGH9j1fbCTf
ADj+ePNG5Dwc1A+iAkBsoJQN1Pni0Q/4Qrx//MZBdz9i1tQRyr8qLGPbtOT0Xuya8f79XLjaYv0R
PrxprnJlsTCjZz0mwZTUPJasoY3ZVnNr47JVKaqaV3jYvaavArCTkIfhczKegprVdUDC+VFReu/n
alRJrptmQ+RJ2aEfPPR48SshLxFETp7ZWwXGlggZL2GHphf+1jF4sZtwRd6T+whf/B8FNakboayX
J67keq9CxKtpCrO71mGhe/GhDetOynOauV9mSPqhMvObKM16aZ/0C5F8Zu7LvY411H/yha2HKGPk
lXivSPwPju2sk2owTedLgdMwjEVKjcwroWFBczbtZkwTM00C4KMQdBBC21Z5pRqN3O6QO8+yD2wX
9hoYRRv0hOk1X8EmC8kKEjpktEJ+SLfTH9mou6zLNpLrYvEu9v63T4JZjs/cUcvcl1RfjZCtcWab
9OvG8MfHxbpg+Qi2XY5OPvfAQE+2gO1uEIePspnkjg0ba6V3RCi87aljqK1/v2GbB/CD536ly+KG
JS9XUMcNJiKXDMwB0Txk+gu3f40vuXJ0K2fIZPqbn5cnRyHnhV/7rgZE//dh2Pp5ZvhtPDTiCCzI
jHV7puDCXVasBdiskq6Hli38FsnmaGYw4kOOOE8Pov3gr/xLpSu6sd2aKrxHYyfonT/lyvwGRqcB
8BRRcR3B4At/2CKEUjksZ/hMm5YQQPaW3e89nxOYJ6FV9xqvacxxxZmY0xrVPG5IlVYbl5ybgQfY
vKDdGYNU0jZftyKQS6BexQuBSvPjSZKQPo7XP9DNVnrmyXPEWFwvJdxx8o8HZSrDemfpXu2WdDe3
gRedwJvkBt2LviB0MWc7RfsD1KmEmi9BrYHahOqQqW5MTaFbTkvrsFrNQSeft7mREI0rjgV+CylS
5AR755x6rMVxhp7N1R8rs3YUwa5WaW3RFOtWApPOohGyD+gb57KBz81sMpa4KkrKyld5EkFn9Lkz
gtZ7JvKBNifuRb4j6WGJyAYH5/icyY0h9yG5JriUMV1NB0orZsoybAcABeKATsWAguLixyXBXF+W
G/wf8WrkBUA6kfPaveFVpoIMsQmD1jhCP3n3K1j2tPyakBEclTSJA+5HW6RHKsZZcqxspYHMhUNc
txcki+UfjYjeX2Ywv4Nw8GQvyRCmXSq216UA6ipHjs3Ew6sUmB5c13Ok8bAccbtQm6FtLDCR5dlD
XpsPXMaDhtVBt+aADFsN8Ke44bJydmZz/wyxMnQCgQD56yLJy2WD78hFlNS6FXBWEYy2MGHCbHNH
zbyHll4ZcNkXNwiF+T6ToSl+QEkbZCWA68eD8aJNBBTAT6WTVGfeefAcjlaCIbqT9/MiL0uy/RZp
Onsfdv3nSE2dUqHE3whe31pb/NNVPS68xmlxPGLWk4yK0Whcyn2xmdg9J6+Bfsoxk3Vub6PnqIbX
umVD4hwy0kcnMjU21w7IkqEuVNb4PWw96kUTqSfqxmmrMHWYUBUdm6j7oj4oBHiJ5Fjx1+HY+Sbn
XDGteK5p54sRGsVMxEfgG6BVd8TAeX0X/1Nu81ygZBSuxEuPaAlZx1Au1e4d/eg8XfXhOrY9hOaq
L7A0r0ttp8Agakqeu8SUYO1vHyIvQvxegqYj68cknLQ0Hrw/tr6SfLPZnVZXby+PtBvPyc8YrK5U
Q/BZRWrITZJVZ2NRVXF2qcOUtAYYuaWEvUwvJejdYkeqkXHTK/BX9DNheAGuaRExtIBCe7ReLg8O
fUrNn7Tc2qqojm3AxMRbuNl7zXBM7N7Ehas6Xq4OSCkmXPM5FxIt6UD/N86DgP3UN0F2eELXGHe1
GtduItHMi1oPOcc7qaxtVLKnY3Zh6Hd5PC7cUXJr9qaL0IOXjDa1eXyxVp/MnnVcEVp5K/xW6Geu
IfgNVe0h5aKJtV7M+3Ta0Ub69zqRKBazEv5v4/xX9uiGbJqA3wmuj5gWA8+MQU5J+tBxKszNK8t5
OfN1UKs/uwG6mFbXMqxoPNuBJUq+zv21/cm73SDqXeodJracNJbMQkYpV4PEvuOG4nrH7weW4B6c
GfCDt5aJnnsBWNixElqLEPTHeiCjx0/ZKKgBGRb+XJwdB5FnZaEeH6/hHl+FQkCz39Q+/q+oiQtq
jnHpwPlyUPQbf14YkOYvHIVOEqwKRuXTT9Dt2Ie48yL8c3lLsgt3iK/xe0qlyl05zNSYBDRMC4jI
/OMu2gQld5KJw82IEeN6Jz4BB2Huq1Qvg1XehgE8heVNrRBjQNzdlpP/A8BQyAMkUKZhsaQ0D/WO
zJ2VzobBXvO1bDafrDkUer3ktPiKVc3H+zEc/IdzL6yC8+LtsKS46QrDhSp8lvR6nc4Nn4+HLlkI
Q/RIN0FXlY0HpBJG9ll1+BCsvXSHe5Fdh9LLcXtYT1Zlneje1nDBKut0RZDoiwJk3bZyTaPur213
hZloCBpwaJpe0a6Fjj/jFpXUOuRfgltZEs/77rxoWlSoayXMIhZhaOrC2BSpvLJgrcoZHXmIzpKh
2GR8qr0kko3I0cCzfmP6JgFpKgivA1jKdOENeqLbd6J7yNJUTb2jeVbpAkCjh3CDwr1pyEvGi2TH
5/HEwWYYHHE51hBqxVS+eryEW5GEpml1FkbHFKDKAsCgRdo1JAwaXysFWUJdcjlgUcbk5c9ne4ht
pWrzVaJVuWX8P6vUr6YhkJaFynaXyfufdGGW2/j2vV+iKSz9ipNeaJ2tSAznrVJ2wljub1FtYZpv
9zr1YegDbdYDZzA8HRP5nQVOvHpVxrJZ6UmhoMKXu/VnjSgHK4+Pc2PZ94n8hH524h+yhCBlxiTZ
uGrcmKJWzUIwjJLUVpQkom71lm+l398FtLtCYQj1cKgUVC2pr7xMiz2UTTb93yfl7wsVPUKuQvll
xNj/02YRogRHY+wyFTEr3mzwpXn0vy4cjwE3C64OQpJxzkeykrUO1d3lLSSE7GBhp/fgDn805AAy
EPsJVGMKlEciwBQySmD2Zbqc3pWYW9ilCiNmcBLKpVVed5+1Jc+J+/xCje+PAFB9gcbXyuay8djg
PCZsXO6NUdgQX2IGqQ6JHl4t9NIP/nfd1nvNwY8L91iFnukt4ry34WcYUdabZARG50N4GUWceGpQ
RbJ7BHJbdTpg/m6JGLd9xc6+FjxnszwQwLSTqjcdIIeSXa3N5nPV4QtOnK6MGjK0bMZqffg747B/
7MAzBhLD7Qr8wnvhMiTg9Zyre+pdCNs7MD1oUfgKNKwgWfog2hWsj3PDxEUyFR8B150eY+F+tQ4k
Jm0aKemaomG2lYT3UWT0L9RPizHiC/rEQROHjjS43ftxCyMIyoRz76MsUdsUswXxshXAXj2khHVR
9DMA6Mg1UTwx5ucA/1Rs0CbGI+9VKlZ4lCJBCFcJuna2gqkFos055Yu1Td2Dzd81DxU7RVoAcDz9
J6MLNrZhvtDjeHT/6/KeCqKz2i3qEF1ARBY/xirBDzcOriP+BMEgqaiFQF/jX4xlCcm4QpdRFm/P
A8ZEW1d57O8wZ61AAhOfS6/LrdUjn7Xz8qzEsR2gDNnech+vDA1GyO9fxryIIyydTo074LDvX72Z
9L2iL3q43bDewivpYWaoLorV1C2I5Y4WdGanKVSK879F2XMnAQr2tB7u94NyMtE4/7JsGiDklR7U
TF+rizvTqV6KZ7YhWOjawnJiu5omCEMHc7OpQAfMLWIbYpk0Fe3L9Vez430eB2B+sNhPuD2NhzlO
EFHQhRcBVZbo6VcByWMYejWptjiGVrNx5MCMfXPeZAX8xZQ9bvlYePzD7hbwai5D4g1j0KikaqEY
sMUGvEZwXO15XW0P0IcqgQPxDCnCU16Uenq/3Kwk9jfubhcDP/WgCgeG2LWEmlNcxGpHQCe8FNEo
oBoYmclKT+EeCSMBnNhmYzlkgdgEC0BOp+0dXO664Gh0uAwGGIHhDZdNTswXC3ibQlyQFFyiD1nT
mGqLMd+DkLXRGUSP3DJ9vl41/3tD6fGga4oEXmlVCglbDuEDjUZNRy0eT6tdV1E5nQmVT1ZWGCgR
9qC4ElbinJEqer7X7RGDXrUrE+XJj1z/f6YGz/InPaYVrZ0L+mNCavZmUWR+LsUzmqL+szbqU0vG
UdgjmyFAi7pGW/KtrZ3eMGl0fg/SCKggeolv9cPw1ZOLcFBh92jM5bs/iMRfpq8wWDt9ABF9b2Ls
fwra4hRkptfzMGkCl4xy7Pc0aYnuSf9PKsuQYutFP0zLkLgg6F+TushbPy0PNy9e6V049gDtOw3M
9nzEuMqivhfguiLZS93v9X2csdV8I+fY7HlwvAb9y7wO2udHwZDKVniQfIVW+NXcocT49lu5HhnR
PybUiZuyeOGVHgQX6gD83TFca2eCiJh3bqGIzm1iATVh1a+pped9+ljFykrUAEY5hH4vkpjYftdN
f6t2e8ASAFUk65bNlfBi7gfwDrquF5Rehei5nqlBZXYqnjs6KcVtPCLOxBLfNxTwH34TbbQnYN7W
a/bHjv+Ac2xdEIVyej+y3vCPCUW4Au5HRlG2UkqB8m8vWBm6xxblWvcO/a1NAu1LJu+QqkGrobl7
IAEDEba+/5RVKtU91onCYqKfKCWpWvkGEycz4X7hzP8nDiOD42HW2FCjtC67Gq0cph7QpLJtq6Ey
nLZmo7/Jw9h2sf2W69PAgdpcllYlhr3qq6w1E0tcJxNCa4IIeuUgZPJ6juwGRCklCYalX2qa1fPB
LGum8Ggn3w0WUlbOeu+z1MXTLrEa2BnSYPDpRNFE+r9hCczyDBseJKaLdOJ297klcCjgoqWF4LOq
MIpa3JYh31r7i4SU+0wpTRxeAkrorB/coyCgiHksGfAZYGeFguzLhT5QeGsnYI7Ws5ITkRL2VELA
ubQjWeRBZa825JmX46EU/9PjGbQeQISMXtqgJ1tNMjMxWn79Zz5Am+ol+6Q1mZdGftEvoTWyxYvw
trYRZA0xnkeGXjqh5AUTlouPEdJ+ztBfOaQNUxk95eOQIUaw/o8/Q6Ajya1UpkKAAc8FASG+MyEP
seIqM8pXCHfIvEnz3e4gwwAlfDQ4mI2Bis5gE7HcTbQ0l+Jp6c2ECjsp9QqX6AWqzxhIPb0e844t
oT88/vU2OYYqOlrsrLvr1MA3rULcJ+k4TJcmcIQKRpTrGWNrHcU5mvKMFzlLPzFbmLTr4rdpc4JK
mqMyyQqyKYJMkSO6RlANre6JOt5kCvTXtJzg+vUfB+mMvO2kdJsIHXCpWTW6L1XFvfkK1j2Vezfw
UKfZM4rXCDwDQw31hA3B9AA8I+eX6kdwMrNOgRoK7eHJEYzX4cXofNFk9rx2HpDPTIK71cWmjgbD
3G6VwnqF4mHlSgu0cBWkEfMv8YQSUXhnqbrA0CmHCJwTsKJXsMpZ32EgNxo85XTUttDErSzHTMC3
EaoIQP2b48Otv9Ruc77GuEkb3HKceZG14aRtVCS6fWrmTGfmx9iBvNN+RxPTtIwBiBrXG0j9SXvP
IoE8Mufoo4BIOaAS/K2ahM8ozBpc/UNKcvsVbLe0EYqXlNOMjUb7Qoq8Vk4QY5BU9hD6AheigBbN
oQIcHQSUuo23+0w0yTm3ofIO52TW+GIta/sKUkOy055ocNcI5Syo9Or9AHLuxsZRg0/6TJsz0Q49
RZZIUBIyex8gBxNCvp1PTF2jpt9/eVdNySfYN6kxofaPDNCzmx0/iMRaMzOgZn5vbXbe62eBm0gg
IrtaHLaf9OHlQ/8PYRjGQQ5jKXAZnAPND0RhSUlpNR+wWJKrZ6+e+4iYXhjz55Pz40lFAJHIeWId
J06LZFzmo+6dwYHQQaHMlesgBZqxwvNqOEEvRQBE+hjdgpkpX+bc7OLMZv+LbzVCovs9opoWAQHf
HPAtgxciycVB+EV1hMMpQ8kgS977ZO+fSuCh+ixUYMJIKQJ6JIuIYamFkvYR379JAkQWtwhoTvxI
gvl2xUxubTxNYmrZb6hFjnePKfLEKB1ZvxC2fawC75OmHPxBoQ5g5JSX6kWcLCdfYYENLU0Y6C25
XuvQAF1cibgTwwFSnD86RNLM7a5tihjkAmSqk1E4h0PeRKTTVcuSGSpapINtzKJpXSJfk2IX2aaw
1SS8+tLOePagF5FthZxVsF8IGE2gb4CzgeQyPbtE4FGk3osd34OqdgTNQqcTi+TMODG/4eey7oii
Tvxa3niHdN4VnJxvczK2gdSF6ZOOf/4g+UiaD3p1ZmTVsiTXr/CZf3wEFx31nIuFymBYkdz6VZWs
bTer8sS3zLklrHhdnLpam6iUK0SBA/PZNuJGMlQLcRyjo1HEmgRC2trg0XI7DdGMq9p1bPLJFu8X
RkZQMgKHMlNR01jlLbyN5akV1JVFWpZwuXZKVFjLynOyTwzjrpRi9+ltn5M/UarryZWWCdMcDG9q
sPz6aj/ovvsfXx9keCx95wW/4uSZ09fk7xDVhdMS/WpvvEmIWKunh+ix8smvzWOqDHXChKd0kXly
BZZ3pEm79VTuzHB/wMsLZ6bDJy3YWJi13bZiBWoZoernoi2TxVVwX3GQq8ijd0BPD3Cyj7eL/TcQ
QnwX2A4YXqw2RK9G0nHiXcakPUZ9mra69gY0TJpqZeDgJTovZvzb4C6J1mFH3u8XnsRjJgDWwzIT
KFgzzXU1s0Dgm9BnlUTz8gGnywXsKauhZKWmBp3Jh4acTnIgscmY4vPo6WS/A1HjrhnNwghdDygT
pQ0WHqvvhfi7miSShJnCgjoCS+DBw1B14HjvXjPP7AK+Dcdc1DWK3EOSknreSs6x5R/RASqHcXGF
kEbMku8gcdyBPq+VuLUO9gg5QKo/E2+BZ2LygejsQziBcOmVwZxDy3eYHdwUetS6WDwxCjgD6WLm
zXVw1aouEXTOaNsj420CXLKiNppzsrKVXkPVnQkraRvC03kz/97JaE4eW1r+lt3kErOYtbFBGYme
2Am8Bmc83k2W7VEWeojJAr3l73vk4UV2WgWn1lb2vYysWSGPuZIipBpo0XU29B/kfkzS0GmQg3kb
cacYPSLLXdTdzKqptj4puhYJyUxRgmqo5GiHSTMVN6JVgc5Xs/ILL4PxTeCrDgobNDRSWKcygzeZ
EaZvxhh6quhnRPDSvnAa+zc0Tl3RD3a+PQrdNnNMRppRKbi4mdDXTHAjV1ZgemJ1lM1XtiTbzSe3
YZNbaR9fg1Trqu+mbPEI39lirWD/PSNaQqYQdeuQGY6jlg+YsohfjrXUqXLzhLkJcsCzkXAKGlkw
FPf3ZK19UPiarm1Y1g2roXhGGfr69T5zxXUp+6D9Xv9ScObExhpNuNcZamCrXfUXmxpX/KLgyIVR
KEjUAhPPD+2cOdFvgsvsl7+7Tdec1740C+ZveYvwxZHvgnL7MhbipVMtWNTyMxS7vnKwekwAhl0L
GTzsoKrwZcMC8+J6b1CHy9OAJU4GZ55tAjXDAzwfP1KtaP9lng9lMwtUxnw/xGQUra865vfkrS2K
t5ZWfd0pdvY9qSlSPwWVYpEOlA9NAPo59oyYkjebPQHdKgbr5jBO0FKcW0CN7VahgpQWNQzuAzbZ
yc1dO25If4CoW+w1+hb9eOGhcUUp+71eSnQcEFsU0BPB64vrKNG4FSa97au8oKuZXI/T3r6jVsFV
g6hPFDM1qMrQiVQXDbIh5E6PhXg8czIPa3Vo2y0XPYzs6T6ll8Rq+RewF54J6gIaPBw9xZ9CQK43
Y16IVt+O2xwy8IlMjfZYDvPoj52tbBHLsACRmSpM/Qp5ChTTVs5kA3xeCLJGgfv3xt5b28CWbNji
FUtcu7LdpLX5V1QDloDFIVuLzhKFys72rvcPWzt07DDZzDdCIfmzLadapTppiybIgBq1GsVWerZT
x2KKsPBzJkk/7JSPoZlaxE6XD+FxYlMfaSuy+vVd2N+ILeno/xDxjszxxj+l0kJ7YSED46sfN1Gz
eojLrrksSAntKivBed5vgbvJLM4CH/E1PR3e0Ck+X+gLfKb8Jqn85faWNrgUj03keG10GU3EL0aN
VCrKefmTob3gOmKBP212Qr92kOnNnRGVO40AwfVwNEje/QfHm0rpo4f6XNSUICieHLlQzXAa4067
1xQj6fmgROYgFV/b8f8rdOGgFJeaF1GcsbFsNKCR/K8m5vsoQE/gxneuFPIB/fARAVHV5UKk6YVu
3JW64XVZcTCMDHmjH4YQmnK97OSpQ+6bwmSCVDWR9eiF0E9tUrNvvV9ZFGjSpVILiqFscsdNpln/
17uWoJ878w5FMkDjb3MtkPklsBeuE7fGkvf6LSgOTRSfu0BmwfmJnpmZSPUyMMmukSiu2wDe6ZUb
T99OexFpF5EbVB022eAnX/lulrWu0TJ95FX/dht2DQXl10TJmGgw48mVJObqam9llaRBcAXzC9k7
sG5eojoScUXhsHTjKhsqZv+q/h8zSdbZWB8QidK35DGD2PWQIkBKrvbmJ92DactNw13FlLInaZyZ
QBLBON0fzNO2e1oJv52c33WAvOU5B1ZA+qHvpdgcbGSJ70guJ3iSvze/NYB6dOkAV10988sCdDhM
lj1ZjDlITFzVy3Mue8sFHgK78QPzWc5C5CLbW70mrxAMehDZr9nX5ukmdObNcRNWo26XzfTR0f/x
iKGCQNdnMEbCSgGwsTv7UOgbNlnL98s2fdIfD3H+vCzEOsLCY6KrZTv3DLxQOtTihgcaJO+rUutO
BLRKJnSEv6/yfBpYDmyOG4Zoxy+VTQYqdVoJQg7Pum9YseS5o0J9U3UaMg/GWZShv/Q8XLQJads3
NFVdhC5GXMyxCNNA9wU6/c9BTPJ9W0tnkz7QBQcQ4zGyNl2eE+/f6csT7rpd39pmlkCb2UNoUIBs
NJpZbRtP/XTmV/X8sr0k3GRh9VxEv2xNBGkRGidDunG3cy05RxxCA3BKi/VXlkguxQx8SNCzpEf2
Mq9GOCACl3J8B8eZJ5+Np4DDmoY3kJKjCVWo6XiPqn1hnqmM5+mqJz+7aRXQiYthTALuOvVBvK4m
ScOw3fWdj0n1oM5TZYv3hat4e4abZqTz/rbA/qkcvD6WIWY7yi5DBcVKaVQKFWoBmYshEW2RWBGF
DubLBFLKNI09jsOdsX64NXcOqxrJ97CwWf0qzWOIHniHMfG++AKDT9J3ZG0VIhe7SsMuSMzb/JjL
GpUWoQv7uu44SZTQiNdUJo+jWlpkb+LEyuDYiqbnX+beVWtCk6zZcLfQi5ymDGOigOZjFli4mrGG
Vtdv1nrRIKooQer2+T1z59wjySR2fyVk5+8LMF9HrrUTfWDI0a6/hqfr3GnbGUgY6C8iydImWHLt
9x928GMuSu9bzd7RCuO3tHurXTfTIDcFfehr4Uv3iwjYgRBlGWZoac1/cvtEMaOWLsV1+KdgxW7A
Ww1UKEjTajZufopzMy3MNgU6jnm9habLLzoaxcrAPOqvB0wkimJEKoY7+uE0O+50o70TfHWOETPD
Sp0pIeRexNpJNJ0UvJjXTBJHpZjMEzhvCvTJTMh1pi91yhZ2Y+fpN5q5AMbe1s+vKxuD/BEp5h+C
k3/gx0XZBCRWs6bd7CJZWYO9Z6a1FbfxGltZyGyo1aPD9/t9AY/leCR3SVhZWTaG0eXLR1gSLY+y
6nmnbh3h2yZT7tc85NDYx+lLJa+65MrElecbQVOyhc7Npcx7gkfABoKK5ZzSnSZR8E7IrxwsyutM
nk2Fmrq00Mc0rYFxQbZqGYMqiOxQoE1KPim/J9gUjbzFOhUZcQRPLtMZmGGNpqman6VKlJQa8Dgy
ORIJ6jtpE3+eBMy7Uk25FyF2+b/93TflhK7GlHE5lgphZmF7oLSIkiurEE4m5ETXNdZ6DSPiEh06
2BUMuLKt1MJj+g/yg54mEiyngv6XpfHvFJvrPEAq5Ay4kI/ZpNFEng/jwROhBp7UwZOpmtuHIHS7
MFEHp3KaGFW0qKOTl1zwK43XTwcsLtaRLlyR3nE2Mx5xhPx6lP6Nwz3MuNvH+nBwlfNKgZqYuTCa
RQq/GF9+n3XJGI0h4mDnHp9E139dbk4CrmWJkTS1QEkRSZEHmp2KHi5qEgMpOn76Wf5qq14KNxaD
NnegwMRA6pWQ0sFSgW3Pjd2g7U7bZhYSaoWZTP8vDCZrCuXDy+QhHWxlHndFRMfLA/McQi4X5Ktk
KdRS6d1ilvNGv2NAUPHq/RUIfhCaZVfQgDfRc0bD/Ixxwf4D1sPQOBGY/m9PeGPHIcVCaUBawPvG
xzonbvJklp4bmNFvEZgf8yn6AcjwRYUcd+hbBRdOzdDSL/LJJkektXHyQf+L9JwA2KrsVtU2v7Ex
1qPFwKUVfwenpimF5KWS56lmMs0ozeVUqfS4QOzei1j5w0wCkzAYU1+iWARULeXgi5DQhjbLCVP+
6RMe7H9efYQ6B0tj5odqLyEnRGhvBCWZ70oanvCEVN4BBX6Kg4EDpA+KATWVpEcSHa5R3gvCcaCB
nhPTB4jJClRJJZ7PoE/90mKJcXmw8EyaSvH4cvcs3xwuPR+CRqC4dUlFwVxHqJYUYY7rL0R9Jk9R
PB5/S7r95WT+Mm8tvwWRxTfxje7WlSbfj23tgTXFXfMoKhn1+kFNzYr05Jsw/oY3UiGNKDSdDsUC
A1RBE1njURPEcyUE/cnfCGj6HiTWDFHb017HZriRiijmIJyQzTBOUABwENzbXJd5NZAKZbQWqF4a
U9BQOAUdPwHrGgDZNV9bPukOiDz+9cIUIu/JhTT/u1OTFkRvQfWZJsf1MMt4gvehgEyn2MDV1i4E
sUvDvS8JaD6XyCyrvFpjVbYElm/nJqPgWOYhN+n6OKE8kB4yGyzCxV53Usm0ko3JjmgRXfe8a0//
EJ385gw7UdL0zEQWf1B9NYfivc0mWg5jTfok3JP8MhIt7VjbYNx3dBfafUL2Z6kKCyrMsjKrDJ+J
z8ygTBEYdgDD2fVAyQ7quQjV+X6XVBhEiORSGOiA7UV3QXfzbFlz35zZycloHqDreF7sTpPGYI47
H3i+PZvaYjZ3VM1YelR/BsDXF7GwkiOVENey3QScC/qidi+BvKBfHsr2t/Q9gyhJQ4Ua+a8BfbzF
8iUmOOOe+RXWBzpMXvlFtBVvVt8sehl+dR5cWtdQZsyF1GPuwQ7355ulcY60AbeS8BlDB0kfhPTT
aIrjp8kMU/0v0/ScEHGolfp27WGXcSngcjBZF3rDTs+cH4dj2sM3onTOClj25IxN8xxe1TzKxvfq
VOaApgin/Pl1gguCrxdOI1oeMGdGk9UiCAkQYLePvr24j7/ieSpuarObTdD+pFFFZrg6BwMOtyIW
CpLtO1bDfiJMAb5DVAST0awaTHmSuzYPQdXMhzSs1ZwSRNgiuMk+kReE95xPIe98lcZNr+DG0Btg
Q/aE3fZJBxlqRHAo55Xhyp4mj/WtCeq85BWbKjnXiq+vD0miICxIfDT7VyW2PuKBwIkXQfJ9I/Ch
21pk9g88GJMJdELEyPjcd9GVX3LKTYXzjfH5RzTRmGhyxEMIaixs69c+I1Vdd4OXNQ1uHfNU7QB3
Drc1UfXSivWCcpUEmbzZv0jFor7UMq6UIA8sSIVckexk7w5XB0LtvrtYvL2cEr/3EthGaX1efXOB
zkWEcd81bEzk5QHI4PORuwWUkk2cwkq3/8qeLnfXomUETy1pDTzyZmQt6lTwBE+32yIprf8m5cjC
gRMGGLESKLlakNVgYiVhQfucauAQhl8pIXPkd8AYqKQiSerxUVrOtbom5BXMCRngWkkDoyki6P7z
ZT47w/hvO4tlraU3EJduFzA64IbD4z/eO+ynKBPKNdQ9pTQysnvenQbStLkPxDg7da/O8BNz3qYe
X+zCsmbmWlD1VmO+PpLleeet1q1dNSlksMXm5mO0WGTSJxQZfWo06kOUd9BOmogFVUqurxDkzX5I
s5PXeGlq/W5FKAboO8bhcl9lZB+suqNKX1wNgoRs/D0kiormsiToZVcp+pSdx3zZizOZvVKj5xns
F93v+Hwm48+9lRchOmAEd+MzhTLHuASaK75grXHG2fk+GLDvDwSXH3KQJyZN6RNqJqWxmgDFKvVb
BcekiXjskehKCHgHwTu7kQybvd8ywoF5PdRapHoFhfnNV3aFj9As9TXCk0s8DEYxdDf2dkEaWho5
1x6SXY9m/oWLb1kXq6H4Ms4TZiEaUsOCBuQ3eW+6sfBrrLZWMg/qRbwU4ar6Bx3GF0RZKrCOGd0r
dg0Nzavssi/oF4TdRvaUapswIOkJrBPjMnGk3Tmcngo8Q3wVnERNO3RdX29DhZ8AfR2OZcpDEhQZ
ItoxmU2DYK7BxJjXPSf2li8uuaUojHuJIcvlt+bTUYJGOOifJG6WuAnKfY9S0XQ+73072vljYxUt
N/dsH19V8+F9FoatNVTBjp/nS2Xbt3p7BwA5RXHtpyJCjUqHAQvNJiirdChD53DX51iCh27Rr/Sn
IlXplz2VNgujl+WVO84yXtozo30ql8sh0dAnCTJzdVm35AWN3L2OdiyipTuxRlwD21PRzqxyZHEx
GYEuqHHWSQjNANl5wjOkQogRbFS+k2KqNpdAoekCFZiDXg+NsP/Ys2gobRH6r+tEpDQ+CiIhk1KF
tXtpzEiZGRw3LNiAeaz2tJUXA/+3RiMbnpwoKtlCKxZx1120Uz5GP+N3oCM9+D4vs8R41JL7Tz8C
DokR2A1DLUOMYo+1asyNj8vb+haEVR8p7GLbV3zcpZiAU2BD8LL0e7vmvBsPEReSbnAec1Wc0m0A
eI/LMFN7Y6bL/UVWrOTL/Bh4G6q7WFx+mxBsROmdLIxRtIE2SrGtNqp2V4gtpx5pCzHkIbbBhojd
S+K+sFGcJ26tqo1hPkkP/3Tuu9EZPaOWXW2OuEtYUgi9l8jJY4J5/Fl/422lDHE+mWeR41T6GwOV
1CdE5W6Z3WjaLqIsM8KGCGAwEn4ClvZsnynaIzN7Vae+GG/t4oC4boKDkRdhe67gnPXd7SXG7tZK
zZOncEzAEaggXrAT1W148iEMgdxLna1FDfcUKwbKi6ZPvDXZynrFDbEGD9BfIoUOie2mgW/i9NCj
G/8L11Qh0J/CrqoL2j04CDvR70QxIoEZVWWtcfsjkiz9ku0HN58KAiRflVtI1aKQAh3CAa0t2VQU
ahK5I1zuDpZ0l6+MgfustevVZtapSnInTwQ1CpGZq3YUAvbOoVTl8/lxH5QB2pE54kGJMypl1lfs
iEYZmDFmUm7/pNr/9ws/DOmCHJl2JhzxaCB4Wk9SAcaNsZuHI9Brw8a5HFMNerPjYz4mczfggHkx
uvwGnklJaU4t/1Ek090wZ8kNg0CLxWbpG/f96MdLNSAh5wpYqHdgHphSM1bBlAL2de+Ik/yH98MT
AOgRfzH2LBuW1I1jBJNUrmjfhSU2Ua8dkhTmPujEWebNN/KIMQtwHTkz9tYp45KDRpTQgCEN//3p
UZNyaUmQkcqNyBZrw80A8oC7xbSnQb/7veHbT8jaYQtLXBx8x1Cj5ybmtfwDJVaTXNyyP61cdHYO
gImHTyFAzu9sx3iipfP8S/fMjLmdd8/zJBbEkjhjb3qN7zV93RRN5DeyOY2KZFjSGDBKqq/vHF1N
wtqy1wDBtui5IDmPxZK7DJn1Mf6LafRVUc5nSDw3mEaOsIGA7IgZsyyyGIDH4Q+9d2ok/B70DAjW
QWSxjm4Yn3WogPhW8MErjEkwXc/U84nMbXpKB+Snd4bWkLFHXT4hqETpCwr4T7q8dFe5nqzsZ9mJ
6DmBvlvzGJ23zrQ9KuQp/AJTbZOrNN8RlVxABhAv4wQogKeCEmlDSrnoL7ZJoL2/gLnfXpW0lRWp
YKlm0gmyWHnXLf4avzFFyocygh+DS3rSc7B3pLBLNH4MYBmbgwwrtbkA/GlOShNN2n3/c232TnKY
B10AnsJSUv9BpkVY6ho+ONHw0TlvqXszzbt2OAzoPuVFvkRk7zbeah0aVLskmz+x31OtngRhrVhK
ARR/6xT+83yeY8NNYsEyCncG2Fd6UNRFTus3tPAoKYVUBt8YhXbC1WBxeIifwY9OP7zRUCnwa1Ra
DxtuxDX11zgBJHJtiU1WcYUwvlGYE6jCfjEM5SbIQIB+8ehFJHfhvoJxvmd5AaiRiUM5Ayvvm1E+
bOCCMLPuLOJxgnSPTr8ft8f13A+ODW3ka8m+VO+1syHOVkyyOREcyE8cgYwIUMKoy1k7XUnUr8B7
xg+vwEi3YBmDZGsRfeunR81oXocvlfONe1Q652puq7/7SO/4rfTwJhOypIifIOzjXryI8GKFCOgI
ecA2sn1r4bketpUXR5dr6gLlR/SEzmjUpC6k4h1wVr3X4P4vo0a9nvEOpkmK37jX6Z2woGvD+6DV
XicSHNaYilJoyiCui6op8/uxZHavUY/C7hge8m94Fqr8Cjz/BKJJQohs2LaKkTQ6BICdV2Nle3tf
x90y1Y4V6KvKIZ9Qrdth8ubP5t5Z6/yg6goOjmZ/eno7EF7rx1EsJrFoY7cDGZUlDhF8fgVaqErZ
vyO8+oNDOE6Nf1fV8/Nvd2dAWSnDbL0lOJKOlNINpdKMWI63ApTHSK72i8WJ7DFD3xwFTd0ygxhq
QPq2OGSesIeRR2SPLjrriTSXdkRxMKzAP18Vx1y8AcZfMMG9P/aRqNMwuYI5rrWi1FhBoSQHUTOh
mxUguC4+W+WeMnkIapuMBM2pkIljnBH9Dbgkr/jtEr4xf2/5curww6Is3O1BB8ouZJFUdzEnBn7q
QO8ipv3jlSDVQsi+sKMvXNuPvmHpjQ5qXl2S95/PeORAnL5z0Lex95/2Fwavo94sy4s7n4RypWWs
x3lESQ64ijBykpif3TmDISkyynLWW1v9ZU3ChOcmsUsXxn6PCJMCa02RUMQrQF8aDqI6XGbF+pwH
nbqoTKoU6b5igSM0XFRs5fStzKx2KzaTMTAqkUCNN3R5BlJJXO1SmB5wkb2zEoMzROQn38STCuQV
Z+PYySdsZqcQHssNs8xIqRDn4RqHhzgy4B+oqtbxv7FiAtpOd99W9KEptVha7FskFqX2nQUkN2qX
IElC/0SyBmIXyLFTYN3Kcp/WMdpy9brKg/FIW//sB1f+10bAk7MXN+tI+CFe6+ku4JRV5sxhiuSL
cMb1bnsSxK317ISRZfyYRqqtaEGaxyuPUPWyedAgU8nlIo6DOWkL9XkGClvjJiSsEeuLi6AX9Asb
i174sPW3b7OJB302b2GEy42yAT2MX01UC8lMORA7E68Khxgxxl52mS3NUxhHR9G1iAPEjQ6B3lLU
A/z+d+ogNxh7Xu+7iJ606QcN8tHBfmh2ZdDowSjWJtAymsEHnd8Ep1G+NUtPH0XVwfmkoX9x/cop
GkkOyrQuhGNkxPbgG3OWMN16mls8TCNLC74mW50rZ89+Kwwxr4OXLLAnK9YKgkodOKDNwMNX9akS
cPykdn1puus8pOkhInQ3XEPvh0WvtuJsItWIp/fcENoJGlleSLGsknkrxq76irBww/WCpemJRUYM
/o7OAa61TJpnCTJdv6knkFjGZ7nxNSrHq8dgSG/6mb6fZAKLtfdJ2AUUM8y30J5Q4jtObnpiOOH1
IhkZG0KWRBiyiXWGmIMJpddilqC0br7xzFuEqRfIpsnKQOKtfRRXg0PX7cVZ5OOureKlh1lgqoOZ
LbzLcYgICZT2z921OgddgU29MAlaJ1QZrxa3TGDGORzRMIULTUEbeNjJd/KPuQvVTGv4d7Xnq607
/Swr9lwImOxCRhgoK57KKjoAZ1XhxVn1kQcJoRInaVtM9rDuEN1KhAow1I7e8k93pB0rf5xAZc86
LD9d7aBu2+sh+gZFN7GUUtBEk1kDhJy3MaAY55HWve2rdLwEzVIFkrRSI++/AG8aaPpOuj36lEMw
gHeli4QbuKoXCaVXrhfnXWffZ52bSpiuoBy+kZtE0GlCwgJizfLiPsoz/zNAih/MVmZK3eLrgyap
0urjEhcKkUgTFd/Rf2JhQcego74YtPjrgW6H8FOxcM3mJAUPGnN8LjlcCvTAitF/uPyjw7o1MqGp
bmgxzB5VhMxNivDNGRqVpd7rjkqTRTTZHw+plabWXpQkLBYOV6awOqjnzUapErvVj9GbC1MP4cgn
3dWXaj14E91jPxBw5r2Xuizh6mkVYhis5NT/R4+BAjzC2prNoZknE6sx5+KBkSFWlTX0fg6VhPfF
UdPFU0NgvkHIH4F1iFKlkwgd/vlX0Vxi/ahYQ0ePq0cI06aYmGq35fZURTf2LjKYOVkVCKHrEgzC
Oo773lXTfIUo3TYZOeRLhSTww4hRWUHF5VmNdTXCYH+bvmrXU6HNK3M9Po1/b/ACis5k4T2Wupyh
THhtPzS6fatlpEBSaRzsY+TzVEcwODIDx5Usy3aIGvlSK0WCrUNwa8Oe94U4D3e2dPnBIrpA5ahf
a6D2SIjwP1kUkg1yV6r5kZditYP4Wpk5XAB2CzJp/UefJvMyy1dd4gvfXtEO0veHXqoIhdvbQC4J
RK3LY2yfRo2xv7P7etmN7iVX/M1g3Jydt1hJFYyeyXjSOneADCvaPiEtUK/OVZccdclEOjedIEqC
WBFDyeAoS9Cj/LNCmiT5Q12IMOYZKyFb/UYkclFlngiV9mkB5SYEpCz7KYpzRKsculnY3uA4YgAt
WrKeXDxUZI6yMxUZCmxBg8UqnJdqKOH6kE/h6OXWRmIuERItFX1p8BW9vYQSkYmszPtulgydFJa6
DlvJuz4libcP704tVUYTMdq0Gj4hIvk3G4iW0UcKN18R90AOYxZks2x8CoQKpz3/iiZ5jfhAamMu
oKJ9BytjYS0sMxZSQTSUXXwFIUWZWb48MkU+ula8e4pubKl5tN5yacU/WwLpTgw7/SEb4iKsTh+j
g5hgV9m0pteT5AzAy4FIfDQv76xtLTiNbCUSr84BLzWwUz0emSEeDy/26yZhlY9n6erA/SQxQ2rL
zl23GQ6D5t4W9kqYX3LQ086IRNvZ3Ns6kZuNmNkK8nkzYxt7PY9m1G3CW/3LJs1HSaGuukPPSxnF
yOi+drzlQKU1Fm6fS+mPAN42bTQ21JSfIaoMzajA8LygCoqqwgkJXJa5QjlJrZwrDXFka3dLzmE8
U7l0pcuKbnjEYjRAmL1qJPdQzw32mtoniBEmhpuZrrpXFn80/MllbtjMC4MQCm2mZaT2ROXHA2QK
ivY2kCH/yt+CII9bEl+9fJQoUoHIKUlj+a3mOxU7C0hM7wkDY37/UiBzemVA8ohoT4XrVqWvhWSx
X1Buo0oK/gt3oeG57wuilQZXOxuRYQubVAHy8DuBnGezX5YVBfietL8rax4Sochd1+gIm7xqi8Hv
8NkhlWUDUDjG5JGF2NL07DtZwyIcfDP3QWbWcaPYHvyP2PntY7rTYGXs8ptM1E0PMtPEHNqf5iOt
G6qjiE+aJwwFPsPX8ezbkGyrYJOU2eabgPmODhz0HgyEE7kJQ9MKhCHPeiZs0x+Y2uY8r04HkTQr
5sHfjyqGcvS2yA9WTbf3++a/79Vy1ik7P3om1eMbrucZ3+FumGP9KzuuxYIq1oLYPvKUJMrXnM66
KMzhxSjxU5xTTuf3aNIqPkU2YXiZNpB8cyPneUZyZxUj88i+d06UiAsRIQ+JMyG8Yt4ro24NYnfR
C2hWozONOgTnwgDxXqMTs5QqFifZ7pjQciBk6KC/Hero2Y+vsgCKnywt8BoivvtMNjTAEj+zXQgC
0Zv5U5ZldTxP903nvLeX6ELTmM+XGExCzp5jAa3+Ngp7LnKpa02BeLrXQlBJ/j+7xoVoDPwKxO27
0Zo+5wDiQK+GrfPqj2od+z9+aeQ0SJ6F2jdyuBCsKaPSz1gRwUHm2vK3y+RPBnX9k+T6o+aSd5Ur
d6sKN+1Tzr5MQoqp3ZKlFHQ6C4y7b6bi9BBx2ytGkLZG7vmFdLAtXQvnunMCR3suNVcyThuLrsyk
lzFunvYkvELuDAhitu6nikCr0+TG+dOdqgppGbbPELM8W+P7Bm4rQjSZFVic9P0lmMsr4UDaryJc
FjOUU20PzGADHLe87MaPSs5L2M7odxJaIIIuZXYtP8+V3PPLiMbhWLdo+pa1KyjeAB8Iqdls387u
YpJgX8x8aJJWZV3SW6+rjqBcVCHm8oRJKmqCv7A0WGWRyUB8dH67A1zqpnGulV5w0/m4l0mZGUP9
Uz8pJjZzhgqw5TfRGpHdh7lQVr/mMwldUbWDToQKSFUCQ61B0YlGbVxFyHljhBnsk8U2jn/2+Hcw
TcOhRP8VZ/kq3e26zWWoLLReUIC4wN4s2IHElGEut2SE5gWmFqZD0Gr/5mylONAabJ0qmA8vVRrM
SJOodoGK5MZVDU3iD/aMQMXuFR/nLpQExnLI9u5f91IxDA3eoyX2wncjlsMIrxL+cXSbRoKj85zq
mfeoj2qWgscvlUe8Xusy+jNPC1hL2b31I2ztOORHkWp+O8buv9WWX36/W3sUQDORGmOe9QryOE6C
wNqRagNsFqDtu00EniwFD9zAtIPcM5pPLc4KS7EHUWbcenYOKgd5rtub+q1BUc21YnoEHJiB2Mk6
c985XRoUMN6AUen8V0p4Xqw0oWNATzGMZSFzpUHYr9gWbFkVf7PxSXb7738dbmulYXbky68x+RmY
/0LT8hTYvp4/S99+tTTl+y8zwcXkVN+bX7/MO0Zi9P1w0lEI+sxjIKhuRalT1eoHF0fEY6XCIxqQ
jKb3q9fRJowe1I2nf5UoCw4deYfuLYU7yQSmTFxUbFLR7bj9kqzx9jUIfTqPuKHswfIeGlZUshS0
+sXUo1mvWynjD2ZshZpv/VcMXeJtuZB+TA9S5HEgsk6mAX8NNQek2hiz3i5a+cFjkVzTG3OO7fh8
qI6wwSyzrgKghGcTirPTtwpkvEnF6mkUzTc8c6dvv+rMZ3W2IKYQoAmKwbUW/GryiF/FA4mbua+3
ylH0a0EIwiEwc4OxhCBhAlNmDaRMKhZzckfWCp6ztrO2f9+N0awwpl9/VtH5IW2LCqkqRDRXR0Aq
NLXibSV7Hp2aLfZYw6/pnDzXpCtVpbbXyAoyu6AUI68X7Gh8fBPLoeUJZUR6jextV5bLT+XS0esq
bVp0UIV5+QN6cqzB4tFgJJsbq+FCVG37pxQlRC+1o021SdaZJ2jMPP1EPatNoC2zA/K63vOTrsJp
ZchBnF6RlfJfpcU05l4VWYplDt5RVIKpC+PClfy3Ba354DthF9LRcQPxpdqeidXNUWv+fqjXtlHX
bcpYq35WWy79cR4ZbYn42Du+MURrFeSPLOFozs/UthFKctV2tORhYseCz+fOS1htFN6Zpy2kDZYZ
QKwRYsbLGIv+x5DlniNsd090JyDgRO/P+xdvjMuIh7MCEZbGKH6TnMZts+i9dxJP1odQ2CN8SnWP
FXyYQy2o5T3q/sUuEKD2rq+lXD759q++rkr740BKud1SSym4IznRd/ccc4vfZZLIYXiJb0bP+1jS
s1TzztqyceWYBW45YLez3JO9BlQ8m/+G7hcnf33hUxOUH27sjCC4pzM5r7M54iYce//FE33ObZNb
yLyHm6MPF6Y20xEjnlfKSzyEKr5LS/olQ55IKRVqqfvZ5a8tM3swHmYPxTqhvKZwSrYUeHwOzZkF
ntvWhxX5ev9ObFyarnxAnVuGvdcOiAyU81RKT875KlM7f3qiAQs/RrkKLhWqd3JNQaQu6HLkc6iB
wOze9/9a2NLzBtYkDpXepbdSDJqpdWybesiGztR7n8ipjFkpwyfZWq/eQz06dkTzhPl2lBA1+IgV
NqHCk+ykH1ftJjxqdssC8xeCgs02Ff80J73yEjEJAG7l31k8BVGNe106tBwL7NwCuOG8hQarl8J+
Sk3zPmB+sX5I//riEMKy0GtXTX7ArEGti5A8DyiA6URSOrwvJYvcPM8KwFQtfcYtKwoEPAzHJ94k
QJuSzUK1fxagi6WeJFJkQNpwdnDHA9gFDU18IAea6ceUbmNXYFHaS1xbvISrvM5qkzS9rvlehDGl
Dl1uU0KzGqTg5o3o9yXtMUSUNUA5Ey0Ke8NQiFTtBp2RlmFHR3/bPLHrNjFvIZ8bs+OncSEWyFfs
D+xGP7CZy1ZIqgIfgb1/S4xSDOWFtBrDWzTQKz6OhJmagIk0Y1Yqgff0QInFSf0KSviSCJJlWQck
PnicBVROHFjQOzlX4jbOEtnu18uQJbVp3yAfDEphtFOLuYiDVgA/fDWzpawDQR8xRDbzciAUMquy
XQ+jjKRDiPbEHrDivM5nlbaKyXbDlHVAYLAzt7+cHRcFMcTDJbOeYrrW30e2+Qv93kSPODpyM0jb
SnrtVY2DMvhkkEZuvj4nGAGw/3i56eRlKF9ltOhLmm3b4g91n+yXGmVC28o9czWJvfeKa/4bMG0E
Js3Qs25qSrKdwKGqdvoJGcZVmm4c/fhUUoUm7MIaFVIiUZRhrb1rXCuVk+8G+1NvEqiCR+aLPINk
37o1jT3gd9F5WL5psaxm/Q65lRQbNVqn9jzaTShg+1EEfdREnVn804kQeaF8TLj3s+595awg2bHX
xWrVGiqJG91vaSClyZKgo2w4TPsN/1cmeGGrsQT7JupyAs+MCo/j/26CAHE5a8ILR2vXgzmecvkI
EWjQFFC2MAhLvaxYqY4eYgPQem+agpFBwM5U4X3DJvT4fOFTEPwDOLE3uOg6B4RnNALmO/2cvl8n
aaLYXcLj/vuiXGJjD2hiGXz2LzGsAHGL4effvvv6RPKkHixVZgf3ZvaT4XE83SOuO15F2gp4CaIY
73eGJjC0fliMEjRuWtfyejzw/z/qxd4/9z3W1PCBIRqV6MayIpCVPOcwuj0fXkd7tueqChJks3th
Q4cIhprRRknnz2VxzDvac83fkyEHR+qnk6uDFSARALhwsyAnZ8qha9avWuXMUpEI8zfEfzXALs5Q
zrTHxhSBYUJMwviLqNB+msjTlS57+ZhgvURf81ziFz1u9fq2jRn1dvl3NIHgMbCQ/kzo8F0dfIcL
NCZwzaZXWmliZpJXdvGgfpTB4fWiVVvD+klLw7xleYnSDJ4yYwJwtS8V9+OVqWYANPNDGYu3ziMG
1J9grZpgGPakK+vG/g4j8whJo5Ttn4VAiAt9uKLFTBu+GpUz733qxJGIbuKjeDBE3IKcC2ESU0Mk
Z8ueltXrmSR2QqxwgGCv9rXCKg4tqBeHV80/xWyj7GTTKs1eWgiKcwelH4Sk7+2NPSpxp8s64oWH
aNDImVrQrZlplIFH2RoZlZ8GBxtgTX2TfUnA0fDgNXooAdp5WAfsLQO4ZvLz29fY40xcncsqchSc
QpktGskKBAZlZOxAAW60O7wpUXoUipvCMJHa9shYX4HoTbv3Fx9/O4zOvO14lGeuxM6/4li1lf+J
XiRDZgHAZeORh/n+XuH2/rxeMKBmsSM8zrIcO4SqwH5tRztFp/mRK3NKj4MMBwxzV3U/NkqsL++G
26wZDUrg7utWD+lPR9u598DEuQac4wsuX93k7cKPfY9pYmaL2VITLGM746X2gr3oFoCx9lEdS5BP
G+UnNHXp44gaFWYPjhPNOPw525uPEnNv0XeZKKt7FE1HrpF+XRnAA+fScSRbahOhj3gLtj+6mX3O
tHLss+mOh6o+u27CUQ+N7Y6tqOlw3WXemionyBye4+Ra2u4VCCXv1RPwr00+bIgq/gNsDWk80APV
mDbNrGjbdzb6bavyyUYLiIhgCg4lTlnwV7EueBaumvjfSSGKq3VU5S4OJ6tR2NAASdED9jRlyvNi
QPMWAaz6aeXmAqnQhDbDMmD7O2NheYpvLhz9V/61TKIpKFP5ME+Gg5Z1SOnXmRGZpcWDP5EE+lVl
XGmimBqq7u+gQdpdZ40mjdZf+xMSo9oH+NcLiA4WuCvCWbZxkbU/cPLUHlmndrvYzKe6f4FjV+4B
V4o3JkC0Mi0F/HS88mAuTqPqJuhhJOj5IQ6W+XNdS2QjO2Ee6HHqnaOgo7/uEzcWmCLvPKNbFZ2J
XI7685P9GI8gD6kqJBlbAK1+/EWChCk4Y+hhHxg20Xbz/riklmUQi/oU8decQcDIxQiego429zHu
K6mqlctyD4wICzmnhzri3K9bY0iE0SkSJDLsPnky04d46iZIczqHpUhiCZgRs7Y5DirjOmBOqyP3
jEKflt/AdG7UR+HY/+x/8P80nTeVv8L7V+tcQLnoVz6fyvAgA6VOgntT41mH2unnOB8PbvPWBLYk
0blnz+bufNeH2DCNEBIcUNWbL0k7F85BueDcCh66RoyEoIbZtreIdt1k0++blHd7+fzs9ojA6tC7
DC1s73b9fSHFndze9kZlw7Q6lCyLP/XLo4ercbU4/lvIOGkx5P+FxJnyvoTjsxadqh5Y9ss+Y2HA
s3T34kmz4vQ8R3EWwGq2Csen3hD5n/uEVZ6n/BvvVJrPkqXlRlcII/bHu9U7FQEfUAxtdgBlENy0
nuuwPw7SLwR0nQGceO31xmI1BcsgLFoLBxBE7SnKsKRhjndTGB8n9rYDPcWXxy0hyVt9lr0n1d8r
Lb6fe9WTVUs2Pbxi5nlPerKc4P3Ufk+oFHEX/1d0b4kIZSjdwmgXxFVcfk5pl9GCsp/kD3Zcjzkg
5QKGGWtuWIKrj9O5xxndWj4S2dlcfbBiEdrFlYCarSmN7vBY8zsau1wfR/nGT/kEntosyOcEe4CM
/q0SN2Uf9DVdH9aCyJ+fCkLhs8t1blS8HWJUzZwcxAqmzKVqpyu83VAOXgNE9PoeeLeZvgAABWZ7
YFuhaZMGpyVjjagWIZ831069NFjWPPRPBOVE43j5PZ1NiHd1InsFskwISTZcVmYREED5JVPVFgtD
2tI+FP7214dA/myGZ15qZlVOkFsT5AP8OnYYH0BbFCfI5eH5U9f6RYsQ8WPNhu28UrRCsa0WA22b
KGs0R/zX5XdWjn13pUEgzA8BMC2uTnR4+xvBzKklR5rbAJ7X7G2zSWFXnt0/cw9iQQo27Sr+CW0r
Wkp7P+O38KxgXbq5woOJtnIyOXq20ESjisVS50HGG5KCKqHNoH2nUVBayDefGNiIjoHgDS/hoooj
L8YxmC7MaEa1UL6jEAqkQYsrv81UfhxdWOt/jGJhqh8CaZNJBAEW8YwSBtkVm5nx9NhMvrPt9ELK
khcl8PrzRNhraM3D9JZUzebnrs7Ry0Yr5XcIHTPspAV8pBzASiBcBumDMEUVVsvkHPJZDrdkuKpE
r9T3x2Zscr6rpl6K38F4opXFgMu9/xx5u31S6hn4vkrV9t1BCVOnPjdMILA8ZuuySxLU1Yg9Idoc
ZMSJofQgCNauI4QcpaMOA2mlbQbiApel52naPq6ZyOo7OSXPhByY+dHdBDqY17g1fPf+gsFdzBfw
Z0pNhKis/VXR71MJGfVJ4kYgDA5kPZBh+kPURjG1Rc0+jF3O6dzHFY2nMbrcug65dWhawxrSvLom
/qIZBbmPcnz444Wuxs1DSrWX87swUaM9MF5zTf+ZxzndncwHyseyiEUIVuWN+UqttJVSp2YnEZmT
/omBaBj2ncNTaFSO71/6Riris4P6MTnCq5V6ZqtH9B32y6WikVXuXxU8jO2tZZS+53/dKaBc5usd
Z01evz6xi9EWfthmuDmEmkc5dAwr/F9e4qdeqoI0RMvWhsZH3Npd47ecZknRttoiVVv3cvEJ3SVs
wiAW1AJ1DKG8Nx49nxUO5g86cJxcKuBexOvmBrGRD3rUcpFLrvN8UugJYEI1C+7mFvPNWetVQEtv
JZjHGCHP0+qMyfmyMjvKoC0NEUY4nqgmOA+8U7jCVT1wM5kPj/SsgMkbl1Dq0sAOTPGoO1IpSkPy
7uLnoM34DSNoMjnU2DOWqe4eKmqauFBs8pIfdibK9hqHrvbAENIcT67GHjOzPgUsOL9gzbX34LhH
fdMD5hunxAvavl8loRe6/cZbDSbBNYZi5vvYj6HgZBsJNPOfECqX+izgUxAVFC5pGW/v06JKWVPI
8R8lphZIK+WQrOiS9bzwZUoAtKvKKaW2kilaAB+fyviIS2M2C+1BuYPE8HXvg8C/0i3t3nMZH9NO
plwc9YYU7mNcXdO5HgP4YriaQzE6QliIzgk2VhB44GajVY20YGzUuLA9D1ABzTndUiK4x3bRSfOw
gT+CWwVKiz9KkORjCR4WovQnLiAMpgoU656HjEPMOMGn5IAcw048BkrIfipQcUATmqGMpuWe1sxZ
/pFCw0ahq9qBPu3pWC+N5rxvbnWi/GxgHfOaFqa1mUHjr4iuvyAhQtykoF5rpBCIVH89DHib2Cw1
KwfnnzVMayVB13u4bATunzsOtkoIsc4WpYUJkVOsSjj4y/pM4kJAjtVFZ6KvMMhNK3Zaq+Vf49ER
gbrMOAQHisH1gwUryz9UzgPhX7YbPkD9NX1EzNe18qvYti4t4nwqVdY/MdMEbzbRNnvWe+NFEr4q
14iK+F7MRL8wwPZaT6uC102Lm4Ix6nucR6Bs6PRGJjFCgB7D7K/n8GmA+9AUhGjoIzsfVgv7JEC4
8XikSTkrW57e2OGtv5NfNmM+krcT/yq8PtEANV8P9LOPh1nNCUcnRUUWfcYIg/WYath1VRWkcqU/
0DN01c+PV5j2TajsRfBvDtqPuhvGBg73buMCbY545/f8K3mUx91xpuVi3GnC5UbG9xSt08KMVUJv
qO/P96K+u3sXNb4vVdc5YboyoXeDRCX4iEBcBc2RYdScENsE4HPagDWeWxTBO+Ctp1SpjJq6SbAj
v8fx342TEOX64bGDoI/fFqgjvZYB939vZEJp7FNXvvOxPcA5lDLqF6sV4clQZuMSasfu87RPJDqa
b958xlSi845ap/MNBFqm1IkC8yRknerMVNkH/XOmRb5PF8XjzbIN5D71GRU6OA/TKPJ4jwbkjgvz
AqN0UIE6hHJQJ3x/l+iUgZhsvX+FdWwuqvb2oQpjHwgoEJvAL/+xMUALyOPa1ZVvzVjhut3+IFBh
e5Kd2ZHkU4wZ+VAI+ufdDxkpjG03O5wNTQuED7DUwwB1wamAC2IYMdZpnXSBWXR1MYT76PBzICNz
j8dxo/UzeudGOLflMbSgyZVtKnV1UCt5CbXRvjbwALdl/75dPOwDfyg8tKrmhJaSmBhq8sEAdHjp
l0wYIkG1wffIrkkgRnPS2riLGTdN78fbsL8aZfeiawAIBTUEfXgHDQKCrduk9YkdtfQ46fTwWNGn
5YvOz2+0hlZfnzFaNnfBW3QivktZ4jlAk1zqLM1rl4R4YqQkUlqlb+lEBkyQHNjpjDYV1FjsNxXE
jvqevYYfGc371jc5KDYpeEn0zP4oFy6U7gVaxGIwkqnW5Q8ZtYP3SnnxU9FNkB1DrogJA9jcH/8U
WaEcYyJwA+xVW8uKUTNjFMIy8X4bycj0Oh7YsigtN1v0UpmwAQ6I/NzszBJ9YVl6Rnqv/WEr5KNp
bviSRt4QFJsvoWcARxilQPN7ss/IELOOdZRYb1fss/ZtMhvOVqKijhGBIzJtL8D2cdO+k7UfdunQ
t/icbBv/UJGvyY6Y3buRQ+S5yB4utG4HgFm3B91cAm//M9VHh/OBkSdZ9tyMbEMnfIVT4TZ+Y5c0
ZCwxrDKAAe0hjn/ieB6/pDDcRqSrao6eQ6yZ3o2LmAfzZ9FF0QjdGTuNrWdDbVnIOl7m7xpcORTD
c4Dg1khzEUGrDbrAjN1UyEsRB9t/kBQ1f/T3lABQOWMB82fQRL07IEfDmp0s03/ccGFPWWb+kcWJ
ofoENOKYHyB9Hj/qjwMLWbporFSKqYZeNjj7fEh9/WWmFpBTzwIEl6vCcZ0wO9aLMrbi9lZPBJhd
4Y3OpZAUZQlZ0E8giJ0mRQDHiM7BEcAU1ixxwpuEQ+TpEvk182bNOiUBNTSRYpe2qBl0Tjgyv+Cu
APFWAZU+ktefbk2aklUe1EomzZXOL5QE8qlskkUtqW/FspUUc1TIk0oBTWEDBnJ3JwcZR14ImyU4
g3g0P78Q6Afvu0G3iVXs+qqXc7jsM16l7TjP9zI96tw49Qrv6cLhnv0nKaqKvBeE7A7/wwItJgUp
8sCWtmv5RJ9Bg93L/v6pUigBFhESNq6haNPB2LLPG+/Q25p/FqfDfwMsSxXXiN/Tffa0fMoASsWX
dYA5dKPNgHVWUTCT+S/H7rMJ45LgYfdzpKp2bigRsmE9mXGAd45ZZnMQ7ooJfP5CIKispYUyhOhd
QHMBWjkbvm7WUUShn36Su9Q9rGkswZOqTYUoEnuQnQMgkldl6dlhNJs5zkjR5pVpz6I2KMVNPy2E
TjDskiMtZ8kynyeYESmwckEQylVWqWPQiftRVQjxCk5S4S/2CFm8vAI+thtluopNPddsvhwurBOv
TdCEB7nBlk0+zvdkGm9Fyh/fe30AuF0wwXm+LD25WHlY94j2gCvR6VNgTz2lNlLVGX3EeXdcxfM3
7EghBQOOwONW0Fw0DYqgrZiptU440SftxGZkEf2L3FzY/gMc2/gIbR2NB982VnxP18RCuAv8yLUw
h3dk0BrepvhSBs2aXiHKp4c9HwblK53DluoES+jcpM2dE3lu8z5JX1cBtsQPPilhsA9/EKeDgJZT
430SznqMrVmWeQZThu+W9vVU8DTn2kChyFsVnJmQbx1Lwb3DPFtukt6pEas2ksjHDIirYC8kZZQd
zmvHOh5HCMjDtgUGZKdg0hwerzaX5K5b/TjMXTpaivtZRiUyvaAX56AbGTA9HRX4EujYyjjE8iOt
M9eZJm+P2j9vKO7PnB/HZrinHGr92DEvt2rEltb80/IMIz14h8vjjZSa9SArsWcbLg4lm5HmnASE
LG2xinUKqLdQCNaEECZ4cH0fFe2AmXh87SkJplWM1kdr1iklA4Yj+PV06TCNtrjRlrGS66nMsGrj
12vLwisoV2vB8+SgS1EPeWIAKAd3J9BkockgX0z5PVh90yhUbsuGcFrbRD2rSXAqPFXEy0DQqez0
GYkTu6YOJwLfyLoDQsVtxDh0Bg11CM9ufnoXcGYSDso8/c2VfF0NSrNDEYZ2Uv1I7M3zJ9R6BYnL
LdZ8vtTb//YChdzyKSreO/56wQsyX73RBHYhIS13NKdb3mvOx1HP+DayuIGh2YZIdtYOup5jfI3P
lE+nE/yAO5hu1m4Tui0j8HCxQtsIpFewwuYgDsx/GzaQU037csL9Rx93JsM7ZGKX/l0dNyEu9b1t
xxcTORxM/6a8h0mHwUJ8uS6GGkaXYUtyWkJVoa2kYeMaI5Eih2Vt33eWkQGwldqVbODAPKL1eA2l
83uAM5L79andf1x9dYuWICw5BUyLqWSq7V7XBfsCcTLDdEp1IKdUORxyBcZv0S4BsThm8E/yV1fj
qkrnAbYw+8mzvOMAm0PWYX/AfeSrkziCUJgQoDpAQwxOnsmGEiHXNqZL0mmT6VxwO3dbSXM/zmKl
hdGMY3E7ouEfcnuak6oVu78X5tk5ues1CYRkn2xVRsF43MxZQtxhEvYlRQ2iqEMgrJLGUBAAu54f
AlWO0Is+Nfrc2TJ6svR4fW72yCEV6OfV3G+d+v0t12SI6YfV92Ndb5JOqfReJKf22kph3gyVdmsi
PTUIjrJ1eVfrhN4gArO3dhscqWKadSnzBzhBZvM4K6IpY0OqOgwzII/82JBZzTvuCn84a5PiFMc5
BYcFqIYfF+h+cDvG1JKwPvZLW6KHAiVAYa6JcncsM999f5y4o5IhKVZBqU9T3RrtzADL9O3J61lI
gJygmiVryM5/hCbaNd5uI4ow0KfWFVBVliPcHSPo9LKKNGzwTwCEYK8tBzTdsEvHWC4oPhbT1tv4
e9xHM0FuLH88H2U2JkxxPBeUIyvXM4mUrgiDwmR8ffvPKjVi8+qa6BcgyEYAbx9nkxqmtdDUWEOT
o0cx70IjcF0bmuR0Exk/48pdfLpkfvCJUpeLNmMr9ekRF+f/++PY4OQyavqM+9abO3KJ0mjie5eb
X28zB3jrYaXxZUs0d/o/8YlpqENqJS4WL7HqU8v+zD+VBo7KYBmYZrEi4pY21oE6NWfHITIAFaVm
sYN+RJopsouBmI7gFrMvnzAlV+UcEdBFp+K0oUQpCTWm6yYcoyxp6tvpk4h9WpeofhC0o4tmF4/2
c2W3h+1FA1PXIhRFwEJbS2jcpr5aAx9Bqfw3C7/gPV3CmKDmvv/IbSdx74Mf5oPrGSII5ljFFtP7
Xy7d2D+8zOTWb9+wJeeYp29m6Jfyvv/moSXXJMUpeSpG/7tlSlkb968f11GMM+2GpfR2kvz0mSIA
xbGbklVJZ3ZTfB7AI2pLp7qJ3wwPLM3mVG8Oy4B7vMIR8RT84qJO8TDAmkWfbwkS9dS0PKKehDjs
WNyIKDNXtXt7n/Ik8gj2p6AP6kwBDUkNJWrC3QzKQAtga5ssfchW4SFd6VHLqT6C0FaXaTXCVyRg
8b6jzxU2D6+8aWHBr75DBM8FkKnBGoJb5w5n1YgDqXtH9CrvHkt1cF0edYKMiI6ktc3or81+Aa6J
gTOZnOcCqOyAy/hgXXDGU/wwE3NOi5SLqUX/Axc23Q+l0MYhr8OspsiGukhiHNO8aa9BkdNfhGd6
6p6WS6aed+VzLjZtdKbcRHOGXBS3hqFkahGB+q8wPNsLOyyN6nisr/uAAx4o5Ftwg0yXOwn0sZ8c
MCfM4un0558LNhdl25ijQBnmqe8BGlFYw+JqRF1eLfY33cqR7TRgjdgs2Kkum0gAgDnbPU9/4L5W
VZdqxwLqRhkjt8invzYhtR83oQdgP9CwCfsLpFY4ciUMiMeH9ggxGRmlBre1Ofxo/avl1o4Rm/Zj
2N7qZgbpfvDHSODppeUH9/rsSge3cAbqgkR5//O+H1S3oBNa4jRTHHwzATEg1oG/6l/IsMWBTRcA
9etoYHOCC0fTnZdtuEoq2nSkQMFnZ7wZGPLy8Np0FMQqx1on9yh1o5EbFEuyNll7mL8sz7FUsIhi
OW2kI79IvFqbfYw7YGOdu03UswfhR0wrqorgB8Fkjnz6n6Ypkl0zKzIoAW5aomdIF37p6OJXiDTI
Cok0Dp12B25mh09dFisk6+GgZmXzh/6FQspquy88DrYlLf+PPFaHgnAk3YGPzYfNyuqOGgsB+eDN
t3+QcBXtc2FfuAzMcuTR86hi13rRGZ3XQZ/qGEAGdX1PviJWhUeeDRVCWQwg4JFo62ewYQfudW+A
nLeM27qUGKG3DFEeWqyO4/bbS0DIVJTabWWbs6CgnvCpNlsxUYjusC1y4gOKVuOnEYiAvYJTP586
OVyPb4LHGLB2j45x298qQuJ0IAxP1IGvKUQFR668M0FNIlePriDH6+QFfkDRjo1MazCwDY7vGCad
olUL1QWVUotfjQy8+0BQjKYWHCLqk9R3jV1QwhWaO7HVsu1OzYPIE7+VHjrCFTSqTLWID9ID071v
fUTsgwTLPC9A7CoOvbC26u9SB8R9wknMB7AHm7Kk01kbtc1COcBSP6cflD57NknKiGEyeOL3RrYL
T3ZV6lirosDBu5RYR1hiqRdIF3RUYFh9h/4XW93FrWibxnCVXMdzrdHn9G7/vUjtEK/ezV6ctT3j
zMod3caWU2LZZrJQMo2/iSVJaVylva5oFx3rVTXsPApwhR0hJv5z8FeaPP9CWN69/TY+pNyKVz+W
1sw6LTsUyXSf5JhtZmAExreHCkDv1nRA5XNb5bD3WwVW2uaeuRF9Nz0sUyVa17oyWiMiVjnYiYtj
bJt7iqgIXo3i48FuICZYXlLKa45e/B8h6bwBXBjlVFbYFWE9pqx7I5Um5dR6fQXyO8m8LgDwUFeR
6mdmZrSGDygKwjZ2M5tgCdhJ0Vj0VSD2rlGuG2+pFv7dPnhHdkyiVpmvBWp2c4vwWXyxt5Tp6/vf
t5Tpz0s8MV+yPtlgVrfcsOnKH9hqPWB1E4IC/SmxxlqHEY0kiykV99h/ODmdxdmiQmXoOxf2D+S9
LuOMKvADhFDCIzwxMLx229mtD00SeAqMjK2xZZVsguB/ld9Pu0w/vrIv6RnAK+C2cuSHUWK3/ic8
XasgdP5z17wVMV0Y66e9NNHDuxpwcc9T+csnG6XdKiEkugPyWPCbb7nQnxNUZiA84ikSbPfm9PB9
aqlyl8Puykw/0WCknziSfiLJsc5zbARihXsmP6isYqyJ3FT+TDUNxSopei/DPYw+l69lAuZfvCN4
nm7jYXymGtshQzmSbYDFaRrSrVFJ/4IDBQUAz1jZHYsLoNlEp34ueIeilzbTmDX83Df72doZugAu
8ChWMYs7jNF948mROxlWIASzsWdbdG70dwUpIc5D9du5q3p0BH2VY7g6zpbw6WuWxDqiAnUuFiMq
Was/oXniOYrVRuUN9XNqDYSknR0/Ld8gvEENzC2tY29BmFc1ho6CKY3CCewAM3UQauqqbQuy+uzF
0AvE4w0+U5RFk+OqyHSg8qLG/BlSkYO66+rUumbt9vxXc077/Ht3HhuETwNMPY14/XqtDsTkilSg
ZdTiKOv2Q0cS7/Agsi0pWKGP9Dva30ZnZWnmZCvd8kS0KhvQkx9YorF1j49jq/PS+Ym/H2CNIDw0
LUgeRHi7yL3k/sPw5BEuUFjsLWlgnoJcIVXRfj4VIirOWc7s/XkowAuqLn1TSQY6pzZImbTQSVjm
3DX4bqmiWf5K5wa9v4XFvkVHmFb5V/TAjm3rYPEsBoJ3yMEHhuoJNbArUMj6ivvxwP1LvkNsuGp9
1CzsBGvJiZiOtssIJDMLGiaZqsCGV+m9cma2xbTGQt3Q6wVLfXlycLMobU3iqJsDhvqNnfQ9Agwz
AmaCuY2FPHlO1zQO13mc/S88YUcnVZgnVrIOwNJLCpnoIlSrWGd+DViQKrOBW3oC97oedSaH7Vm0
ElwSkV5nhnER46E/ESdJ/2GIOqSKUIhFIBv+9YuVZJjUpocxBAEhm3MpgEPWuFPUarF7SHzSLuAX
4gB5wTEJaDH4d5mabJaEIhkQSDsy1HzMRpQ5++52jHdvd8NLp7/W9s3cru34l1zcOUFLmS+iDad7
5N03ySBHFrwg5Aj68AKVR9nep98Gcfq/vIzwJeV8IKnTL9k7TiPuKG7es5fFzmvLincWMm9foYd0
jAZ9MLWbM2q87aGWDzvn1ePiZa18gn7gftLIUkysNCM4zrnIkKhRKXF/g2p0u5c3vOo2zTQw6l9j
ZDXXFb0G7hf8DFuQPlR9q+8hidIHCOM+tweYx5gvqOQiL0YKw0tY+q9pfbA/Yv8fRkqNrs+wENoT
ClAvIyZdIwA0vVZM2LLiVf7SGUoewdNVn1SIG5czg0Dxyxj6CDv/mdMw5c5yZNli+HOC41MnVH+7
eRdSkP11beW2gLR5gCPcl3/SzlXAeCmauAyyfos/E2WrTG2aDYyO3gSDVrNHYpzWmodA3lsvyPeF
hng6GyhstLyyuRxvnaxiHY6IzOanUcfzRnQUorFniGtEWn6gYWtbJ827BD/i6d7Zxwhvtyy8E6mP
OGiDw0NtibtseIb8WtTdXZUd1sAASg5TBmuXZmgStp01+/oaoVI8fFwWXwehjJ3k5+AePvJtAh0g
eDfX5rHcZreYXe4f19WU04NjnW+A/GSMOIQFXQVUYDPFhwn7HogQv7yn9R5uTzQaz10TG07DpbSb
wEjjKsUvkXAn/fkAQk3sYQgzDYia/+K1A7Y3QGi2b8geiI1nb6TEUsTtAIMjp8X+ZNR0246v6s2Q
bJ3wTyqE7upgFa9xbeioYFlNvz5m4XjX3QJ+FG7eS4CxYqPhwmN4gGUSVJL5n1IHQEkq5XJkAm2w
W+6w9aTGwzqTAAPN0QXQzLf0JfmypSNp/sxow9srpcGuvxEuy5TDEuG8IAcYjhVpupEjaziDmUNV
pjXBqIJE5CVx/Z+wpsGiSfewYLUNeLwMqsfK2JYLksF0irhXKqCmxRjWxGUqifV6RMl5dWsSIAT3
tfnW5+bY+vRwBKRvvJNczizT/t2B6m8/r1n0Qxm4hZZSMtdVP34nhTPypysDVqo9280YxicHT71R
uAhQJ1zONTXFTyptNq8R6sXoXrxwy4WIvpp0BOJnME2ommz0FX7PM+n+mWKG3ISUVHl3G0hsKPp0
L5TY0l5ThToCTyY+OK7Sxd/mYNnYlhfMAOF6YrmyS6VDI2nD1/5b5FrOIJtWLFR0dDzVYXbUn30Q
r2BYoRlVIiZFtgkd8cpu1mR56wv+xG+18WhgKYegn1u/UZ9ThC0JS7M4U0fSEjC5Y3HKOhWHe1xs
TF8D1Cb2KBKa6Gwd/DDg87EFaq1oI6dqm3Xo/2Vf+vWV/f5Kq9EmCFLlKUVoUoqqWsjqwo3m/C6o
x/yLP22knZU7n6eRPKOAh56X/PHSAn8RAnpR14oAftwJJDCZnLgyHlpoMSeeUGwqX8A5viwFWCt9
BkgWSqKr0xnFAsuZhqteVmN/dKPy/C+ybDKygNhK7oeHWirg1xltMKRMyRMzZgbb2joXeBxFNNES
2DCO7g8zwhcT6/h9A6VsldWpjQ/VZr45G1rvJepDQ01n2lSQrzA+2SNJb5IrjLMHY0OviBDzTnH2
cuLotiMGrdLOlw6bYr3Qp6FxYNXm4GfXTMnHwlh2+h95BMl0O52mMcjdf0DG6jx53gOCIRzxF/+2
402RqK+uzSTM9a8AuMNOqG6NnQm3jDmL0H3b/tosgZH4kVaFN2VJwLXtMGhiD6TfnQiyQZ3GByYq
xOhpiymLi/d9+urND7RgxvUQPKTfZ+E4qWNWDBwjM/CmXM/dusAGK6WfRabm5ndR10pgrIsej9Ml
jsh6c8E3A35lZWzKskLXiwOkc489j5hcJeFGqRXsuRRiWOx7OI1R3cW+qiP6x45CLI/6mlXOImeC
0r936CY+DiOzGYusUFGuv1+2p+CREXNK8HX5mCy1vLmihk1oJ8jXQ7TNnYV42bppv2RvfLhU0P7G
f2hl3ECe1dR3euUb9eqEA364Cv8fHbl+ou4WVsYoOxlhZEXXIAPd62QmlcanBwdWtYBCYeOHcpZk
qYB7Ghu/44wiGNRn1ATHHcsdS/qKYoenM9ASSzG7qoDMyQLquP7DOLiYuZV5AlYQkoeLY2/DxZau
W0AGyTw6Lqtqc4cJZP4IT1IKJlKyeZd/09LNfFOXyz/ijgURy87CIdo3FNuvSW38vzmeNy/6mZ27
0AfeK2Go9eIJKRU8If0PWTA3MK7JA/Lmnm1jFMn9jO7NUhP8c/Gd4t8jAggiJHQhvNOuNpxCypWh
lEASGo+pOHc/UAM8yO7Snm/4oPadZOpDboDi51BShUiBXYLlLmoKmOsjR1BC+13qNcEXicRn4AZc
koTFqWCoAglM/WOC1rgaksUMdK/DliapFbl85uY8vcvyO7EOc5Jp5N7Q/tdjkzLlfPYCUNPhDVxv
w9RjPX6nCNNg9nlQd57JRKebk5JyWNXTz3wIsgFryS4sqYsKQq67yHglyytzXarOJ2oFM8jb5MCs
F/p55snf1u0l+myDrX0EYYWVDW9lRAULrJ2sYg61/SHU+0UX3uwaNFjlHeG2K3el7CzcXgJ8fnvI
QexAf+OXW+CrHLOwyv0qhzcmkEVdLvU90NTG/mdFfoOiSMYldjfkv7m9xQmIvn6Kqafjx1Op6ePs
gTKZyOGWCQ8ltQqE3+210eg17lsLFMbt0qcrFF3Mw1WXHVtQ3fC3K/G0J9WxikQPFcGbWSNdWI18
RFVMtiSlU9dpqquNEMBPv34lkGYBeaTL75eOWjLBVm5Z+oMvz5omUDFqzTdQfDlwwoijdGRJ5K0f
nBVTZa1Ge4azDDL3FHI4G/lYHCKIHNVIft1HSrr0NWU/xhagIvnygmKQVNhaIZIz5OBoQfSRatF3
xEOKir2Rwaf5bUHCMaIlqNI9YWxK45orbG+U0JFRwSXHvEgg5Qbt496iQ1Si3u+LXd3znZ0iNwP+
llvYk8BmozvTbP74OHY1G9mpKuJJU5UiwVhC+tAuzd4wMj3zz8eM7Tjyx7LjhwU3tlxJSVMDIXev
tDU1WrGDKKiBQzpJKAyuZTYGWF8vJ8Loq4DQxwLSlKaBFAaDhsoVJxlkugMgt7e38sbIQsg+0f+u
KmjO1Dsd70VeOF37Aus+zBuL18PXphLQ703U5N54qFYzo65gJDOQj+1cj1jtbjy9PR8xGzkVyXRG
Bh6zwj3+iiPG1XWbU/RxnwfzlpNVoM40LvgfFIDKd2wTrFjRokbDhLZpG5vH7ObB/CFmSPOTiLTQ
2s2i/1O0N5VaoFXyRLWnfGn6BT9ZDRenFwWtc/CzJs5nqP5dS8S4W1tPLAxysCqc1xzQVePrkJbn
mqt3IcTrKJntLbNRvbHelghf7q4vAgVJls4oR1o2d1pyITzEcRQ+Kxfv3NAJrnuH0cRX50bk86sJ
KvWz/+iQ0wDZD+gNdUHvgTsJfCoV+JVkUhO5H5Iwef5+QdpmJW2NzMauD71VvQMfDbQXhj8yuv4G
jsq3I9T2WhEy8TYIPZVXo7302W8rZyJwDm+V54rJgA0lPneEfdhauNhYfVl7Dfd9TN4pbn34xo+5
avVJQArKXnDSwpdGAia/upoZ2oMHendytBz6djepvNZYGOQ7EQ56mHoGyJy3ggp0jtYmAVvkKdsZ
KWMHBWUYuz6vwehUw8FKl6M2MT0h6i5p8Dhid3q2h4qRHcOvmOqsWE+2dYfg9oZ3sZQ8Dein7+3w
aUdv4jkiHX72wpYuL3P25GeC71MmvsEONW5Cet59ztGqfE0MO1aTx/sjfYkkgRFgvbZpnYyhqWq4
e9Jv1YsZWmvhDoIt+bOGJheaIgd/GZ0JgcZ+hxDJahLgh2LJJcXdMlacfjgsjSVSb5dY0hSM/9+o
h/vni7wqZvU2GlLd+VttEXN2txCc5QBqPi9m23firB/FebavXx77lGbYfn3srxyg4bk3SPUwnf7D
VP4s1bonBESdFWNuMONqv+bstPYKWUAXOC0YbvS90bK018bJN4+s/XwsbKKlRN8hqYKsyBWma3HX
EXfYW5Ykna1VJAiqP0g491Yl5fUZ51NEJzJmOK/9fO0IY7TwUYl3YNG+gIIRiAq5eaa05YTLbIbK
KF3d5ivFeQHshLM2gRGxoWEcEDNCNgqYwjVMl/4JyzpGBJxYYCFRamEhA5E+veBfWh711HyD+C1H
UsA4bSdF4Eeb78tnpXq6+lnrFYp154jaB6pOzPABNxbCM3+WZafV8YVZRIOvPddL4PNl7invsRNf
h5HzEBr6xI31rMQt6xN8z/FU7lMsT/u8ZulV6b0tZY/M6bu8IHkGlZ010sEtt2AROm59907DCfjl
X9+C7dG5fMoJxsXOoVGJVrXKnjCSVNKbephLNu0bHCdlTbbLcrv7tPK9XpkPDpNpRmnd1+CZr/vH
C5++aPDrK9bwiVblWDxlLuqLbUcvMHHpezMG3UMkPg1kSDhj6lavtRdDW9igm+Q7TpEqozvzf9TD
vNtBbOY6XuXOPlrgEs9eLOSwCWoqM2RTNfEFx2UR6+1j75w33sjk79K4VhEjtu8pHHgpmGvQ3ljL
yUefgVFHSHBfB2dMUsm3lH3rYg/awUGZnEzSfY2wgEY0RC6omihoztsNJuRG4KpldKhUsEUK3VLM
YhdztbIPBMgHM9PqtePoHqhouqcSFwHAaex8cO7Xmb1N4vBlMfHaa2VGFGU0Ec1l/r/8KnMEEjZc
mU2S3nlXalcaGSnGARMDNj/kBiY85x56iprMApKSpLExtvH2tuAvcckMpXTosXMtWAlKo9BTHeNR
zYtLVF7+IoTv8LdLGonDv1dpCQPBOCvgqGSJ1P/G0IMafQEVzav2xONPe41EHgG7jYaERHQrjmHv
nd+Yfmn3INgigO5JpYqOisJLtEuhrps6ONBSsq/O93ETOHNymLu8EvpUMlyaUENb3Pau8mgiXDY5
C5N5AptHvYtxbW/Fv/7Ttwr1jqOXSLtVaslthTZPP6FvRW/hjWWXrd0oAvjIs4vQyKENrSx9WCkt
6uZSZtdIbxPQS7muYPjaHLg+tohmd4dGwCUfOepp0zNzzMQa4SO4utrTDSFFaz8zREExwqigk8+w
utILuWlfBAtv8NuiY4NM83umki3B/UKC1Bu9eIs7vUjRm5gmyt/TMQszU2yZB+yugk6zi5luhjxW
Dc81PYfFNbZrxItT3Sxj/1CgM4ggSrx/gV0GCC8E8u4AfJ5sD62KBTSESTBeBvCwO3IYZRC5Z55i
iYs+lS24HfSadVvnoPqBHFbl6aXK0tXas4QDq5FnOhTwtMxYhMbjqbsa9HQ0Nq+fzh0Y8ttjVc4U
yYXEjokAqWSoV7X92MKZ1Krv1g84FECLZrf0QcAupjD5GvJH3rkxB+WaYn968M3L6IYaDunlo6Q+
HTJ8/a4An88MosEdSai/MlRenbz0q2/CS/E0R47i/4lZYiAnLi7DL9OuiYC4TFfqp2tk4F4j4vFY
W+oHIotrOInxu2Cj4aaDyht165q/ojixy/lWapHi3f6QNxZw0bJkJBqYE167YhP01iF82M0pj19q
3BDO8hJ5xRwAnRnYSS9t9Rh5w4NvcZBVuamd6R+IK88SeUUF3ghkL8IhlYA2IcgcoLmL9Ck/skmB
O12SHOIZFCRe51IhAah9IFfi6xwmO/7Fk+Y/HBJUaBH2vyo4lrMSZXWnzmqjMD1XMBoxCdvluc8x
DPBxTZRXauWrBYkrcZVFGz7GMm5yfIEGhpRbk/QKUp82jB6qcp8Bq443YH6tC5dtR/uSzkFVMiIZ
9BoyzBcb2k/X5cRLT3ectIyIJZXpud3hsuYN6rW02Xtyp4tPNswjWZhsh18d9T32dDwSo4k43k9v
7yRaPQT+qkUFS3Nl0aPjKxAjKhGcEr+ow6B90OBZKhAj9CLp9HA2mrFMUsWgVTK4nN3ktlParCu5
rIEI6DUDwSPi93Fp6ca0U3dcNTmZOjcCN74dD+dE2ltgr2ZBYggqU3HG9hJHOxgxqhSl7awxeCwy
AflnOBBb1+hyZ9OIFGF9hPRd30oDGWs2SedOR5jZhUNe6R9Q1W1B88fcKIDBLa+JmXWRbVKOczjm
d7FAh5ktv2OB34JRhIl1SRx+SJT+IhUxjNKoDu889NrmwK/0Iq1bt3iPN0qoUX2zlyF/VEWRa3j4
i0VIXnOAgnyEe99RSQmu/o0C7P4bn5wK6A04so2/RS1qrf8BYNhFlKg+aaT7RY7tU7qR+FplWG5V
NvtPNfqVFpDYPuU3tmSomhqFVr70BfAEySsXqGlfsLd8aWCjh+ssYXPxCkUxqHIBq7C7uzJmWaKG
hu8uXO+oc72kEpwvewZjwhr0A4qXrhKw7CezxwRvLEXgqGZbYsAGL0OtFIo6dE2ewzenpvTQfqTQ
cBfdYusuc9k8HC6SY4/XybmGGWFX7J3Y7K+he5L9OJfWcRox/e/rXJr1d6Ot4elqlaM5176AffQz
SPVDJu2739iieu6lcP/5eH5Ejf61y3i1XHXSkJpb8wmIrrQk0HQiAVMBsIJtiTK38U3SZb98O/he
ikE1mPdXKZvBqCp1Ytuc+tk1NNIBmxvjejkrrxQQZ1WuNir/xEIgQB3nxoHYnIiiiIBlVV8IBnSr
vahimkZr/TGjTjXH8FGeZAb2F3wP4Jn6z3aKNKD7TKuA+xtCKvN1/hSD9/ErfXRU+lunFDMc1Alw
dhKsX2r7xQl8fIQhCE5Lmx1fl1WxHC54D4cOkVYHr8EKcRyfUkp32YP9/Rv8PszvaPmIBMd/TLtS
YG6YXRegjCoVYuMPf+Iz0lRJj77l0OllmiYj+EjmNAcqBOGv9P++w58oGrgHBZfaZqMHmDWAp0fI
M2iwdTzP6KEyiTvmXP5rSVP9LRgGa849238SdNJEb8ObTaYbvMs+1Lu5JX58BY6jgIDh6o+0viiR
6PJ66v1eXhHHZPX3nrc0HO43YHLaV1D0aR4tyznV4TQn/eUFbFoeGtodlyyxNyRWgC9jxUcrbqKv
zuPyYjiRLvwJjXudiN3pNzyQ409HUhHjQ/Icei02rGheJqansaQziR1R5jAar1zSUBqFyCoi2eSD
v4ncdI9Af6ODZAU3hrdLDGZugkmkTx+487cmx2DJrAOjYNHsKyT6koXI1z00q9L/c+vdCO/lsJtH
2srC5l+aHruezX7SUzL9C1vGcfv6Sirh0ufvfqivRTTPeRCxBOio67JkYbJhko12pl8HHvruSEJb
v8v15czWxZTpQ+bJgr0auf06+xJJg4uO+hOLZx9IYvZHttvT34jD3IsWrH6crVogKfztMivR+X+H
1kBswLLHYJWzHA39O+chUS72zHuWkGbp99XMZnltGsPFJMIIAZI0EIto/cbL8ph0o0o8YzGJ+JC3
nw0QjaQIBkit6qHby4mmpAu436ILR16eZiS1j1f6odgvYIJRK4Q76knv9m7Ofm4eTWSYO5At5k4g
CjtF9WQTTNM7pf+pw8IeMaKpn1/IyPBp2Ql3e4mOkVk+tfx7qSpN1IHTIKQZMxsfuhr7lqbKYc26
gXPD7l7BpDATjrPGjgKauZ9KVRYkpfGQXfl4FXwYpxx2fvq5fJ6V80H5U+CwnZsCKIyZBrnNavhw
vOvuU6ENNsAf/3PpOIiIAaq0ToRNVTdg8Ur1YoWXRW0+7/tP0FN9xse/MWG3qOPJxenXKlcpeSwp
J/GutkLsIrgUZaPwXSdZVmvd0teVEUcwWdwZwO995MBlqmGE9ahRJzLgjQngLvEe7926/60QZYB6
lBxAhkje6qsDcR4s1D77oCVOIMJBxOZfDQoZCUYM4RgSUk3BbC8wLV1n8nm7XEtkHlcNMNOaHlMD
WwShpUwabDC5E7wQ796ya1c5hY+T7DzPBscsnzXVX1+okeQka2v/0c49tf1JulwNGUoAFfimQ2pf
fhI++r7GYdlRk9cgOQiVMhGOU4cMDk5Nkyr13yAGdubkdmrzU6onryUAoYoe0NIPfbo0nUo1Xelp
/EltoFKjVoEL9aX5k+j57C5bl59TVlm8rlZeMCSuBDpEXSbEUH4uq7mWigJKC6hIfaAr9Goov1Pn
UYay6WzxqQSjs5yLpLkm4IFz90hns9iqJjdg1lum6Y1dRBT2CgtNxW+cYFCamoRgflzmrgAEVS3k
+1f3+5F6+WNvyw7zbUnEu9P1oX3ubELJ4mUFAER2RzCd32mOhJLq+qOruWMFCWYiU+0Bw2tfamB4
uT4AHh/IDf528fFYZVmyiRPIxHMj6YrKxU5ZsgCiL6umtQnxQYruBmnTqJOu1zDhHC4c80kl/HZF
M/hNR3rhzGiTSr4vxMQSNTsExtLBATeZhnjVhFdJwkXEX8mSLz4b9lefmf/0B3naT3CpiJiBH58t
TV1BcgjLLhAgQSfHwHJhmh2Siwory/0FcgP4GJ/paRt7wKXAFmKovgkN1Q05ciDyp1YZjYx233cf
aoTQeUVE2E2DHP/GgA/UHoFciW5IeE+hM2EUFk8T5V5TXu4PbsOdYZtwaxA7HV7iW6hLa0ttowdZ
P5MPBbqUAREH5gUq/h5bWL6LELUsNgUtpD4iO3xFIWqZM1xntBHHNC1WTdI1scBuVLxQpYwtSfpu
mvfa5MSztkC54kzDYrCqVvE8lBYKYAZFhtc5wzqwpYVG2o7e4qpSXMhZh9gnt4OO25+wHOtpMnnr
jklR/2fSIb/qOJagU7hC2aTS5P4r8g2QLkdKy3TRNe9YmvmqCibZFMt9mZW8gJWCwILVfuIcsMDy
UBWamtHsIgZ+30C3rg0PEgows+h9oj6s0AefsNYcsvfkBtQg4zdj9hXw+QBlxQhWU45MRJ6Oi3Ez
ad85oILsgrdqZ9RqyoJWfl+luw0NwbYaoBeO4Om2XRBrGoXPSy2PcOIEbCKEGxu3Pg22JRD8TBou
8HOMh60l+eiLZH+FVF8hAG0x6kvzDUJosNdYLVIWwWvzVYoTtejRPl+6eZGtHlfH36xwkAO6CVJf
9AVdY9oaTPa33CVtMPktigE+2/XI+hal6D/wIutpd/47OU3Lo2kDs24eh743sQqoCwZnvj8fA5Mz
bZk4BA5bxmoT7dCzcbX3TMe/+4NTr0v6SWfCIa+P9PnMPKS8hXqspgpo92A4D1FU6+prTJQT7CJc
VVefGs4wBryAXXbeT9YlEI5CsgVFlwhwtb79IxED/DmL81QNWodNcs9geb8nh7rybcnfrE2rMI0r
CD/kr+18VttBxtWMSlB35kXr2Xb30B0+x6P1DvOhehuJLspZHfthx7g27Xs5oP1mrNm4loTgK6/s
yxO1wHBzcMz3tfxP9cpwiQrJIWCv5IBsSBG/XT7KoIl6vb/tf+yuJnHROvDBz0ZHLkktAEEJcFoO
7h/KRnzIrj6BlStcJWKNo/gKssswA8xGAC5kOZuErnQjLzslPM1wfits8H+utskbQ7KJdABufs8k
gbtk1Q+61C+qrcPIzd5LAQq0pPrN8tsaovd+ah04u9/O1b5EeDpjYfLSsFzbIs0i5dHUS7JiSF43
OKXy7a+XTSeWHDPlj94ngsQgIFgnxRInaG3EwpMXPOn2lv+7xd2/czvsL1IfulvBfqdH3sLK6RQ8
mipAkvDJHNjOgPuS4oacTM9ptpzpwC7EfSzxZIKdZkTCj+MSF/N1eMuxzoEJl3Y6QaS3umUDz5WG
eo1BCBgifBx6Pg9EM//NjIPNKE36dkvwBWoGDFGIgB029luw58JUR5ukKFkAq7Ccdu+AHXhcTI2V
fL34tMOtO1K6WopYmgSRjLddO+D1QOCIUJkII4UZm2Bs6RqVKqjo7pltisvyFAIq/QgQbGZiERxx
J4U5njW/uN6Ul5MsLuKNqkxd06stffeaUDp7vzUUouWQQ/wE3SsBBxHmeCFvnMk0EWnrkoy3a7FQ
XvNJCGh/Ft7MaPwaH+D/AeyWQBysof4y0dH77WidYmRBLKgpM0a/mCpqzX7o6mEYIXH8cjb1wDwX
iudLzQKr1waubucUknrBEnyomZO5HwvOSgHnLRLYB/HqdTeHXqhKNq85O3XJXlsxkmkh+M8QMOmp
m+B1ekPRYX2ra29LrWHJjt0Xz7kNXk9yXoH5H0m57a+O1REBOJC4+ym2v+T6CNlTZVfsJ5DcnCRs
XJG3K5oYP58b6ba6ucOsTTleDf+13C0aoCdEpFDf9SPj/ehAbNHMucLD/RCcP7knnZpNN/sm9XGr
qeaXIzO7RuxYT/YQEp+p9UANJBu0W6VEM6Gn0yQaPFgd0Hv+Ydjj//CYYVX+tb+c5kNl5NjaLVuY
Zxw3KMC92y8W1ZPyrpXDTcqWo11vayS0pNBsdTwdejVz8NjQFAEKoXiKmJhSBJXE9iKyPsj7trzl
F8EveQxDdxenVHXGc4L6OuTJrYq7Gh1zNgpnTcCD4bC2/iPpBg6dBCLyUVzz/PICfg/T2D2GmqA0
t7BJ8VyH57efx4nr/gpT3s6KaT7tSHsxZ6zrjQ+DQR6q3vBjvSEm/fwuuTq5p3UX0SvCUo6sF3pn
pz5mbC2qtVZJJqva4sgjv80+IQj+6Y7BIcVFdsMAGgfdXEfULyqLTKyqGIjI0Cpixj2ye85wE/tb
Emr2+0xxonEKVOmJ9UzsmBoH91NLD/9a30dpoojFT6L/JwpEVMLwAdKtPj0wwg8CmUOqkTwRm5AU
y33H4I0lN6l4+tMpG6gZXz1NKpyqB3vwZgUsym5sDc02p32X3Lc5S28EofT6yLPSFjzqBiptRMjz
pabIXEo+Jdl6WtbZUuexVBaMKLR9mei2XYTmWvkvxeU+R+9FvjE/UEBmSq3tN8hPi8wV/lmtrK0U
6E9UfNfs4cEQYxpvscPfJ1eaQ+ECJLDmmBLyeUtafoxlsfpX9GSovcqFKoVQB24YDyvnkD7cYV1k
xzNCt1QpZdSijui+WsPgjRaWTTXNr5w4EchB6QTOj685KdMVwX8uhbSFCERx0DHhkFOmKU2dePZc
JGV5I6YsBcrRcrTJPkBvaRI0W2YE6t+2nZPPtaxzQSYuK+Fk68evD5AKN7OU5d/i9O+DZ1SsZ9tl
eAmuS0emsc4+2nop61b/uu3bMkfI9w37h27mJzkZeJsD6+uHJ1mIkv+wbZJf0IL6CJBXs4iWvBZD
p9p5fYx5BcZE4UQO5BVpSZlQ7URl4VLS5uDVI4g+wAxfQ3kqD6kvRc/FSECg5mTMTMUZs+Y1klsO
qTpb2mbyawEvkf3jtXOg+Qq7mM+lEykeimWows+BwiKpCwoDRTENC5UH7hmkQPkwO9s+VJKTfYJ3
pABYuu4DdK6/qsSAXLsJwTANpomZ6V1HqkHQM9r64L9tuLxD9g/2PAT94IxfBK4pha4EKBnzmzpC
sUQ32WQKFJv6uHnyaeXDC8Yro7OjtyXdR5aR4Vc8bo0YAy0QO9eKY17RFqYq+tRwBUeyRTdmCYLE
Z/oEUy1SnnTDopYFilDtKb19UP+6kbOGcLP7Eq7TdyCyJzE9S9PElvEKgu+HIAjxLBJRIXRGovu3
SLyWDPUaux2ZwPuxBrgDOukzuiM4ybLzkYyS9y7X5BcDDhVCIaTv2HP8grP4NPwd8ZnUayJPDZSE
KBCVdKaakQfum079iMNH4guLweMRqrTZK6iWK+DVjq2+tCs29VEdy5pAtDF1NZIHxuwe0QNGMnjR
fn2mvCszUFuxMbVE2ZgQ8DAgVmqKYFtmX/RfGnODst19IFCFL04LE4ctJFXJh34LD0p3zsX0uIUq
SSy4ndPFJyjbRFQ2ZrYyUG/EUHnYg+XKohgyK5K4//Y7df1IA1BkV7V3BUu0KA7h4T4dcFSRJRur
gvpJzF00brizWaHZBFvisN4Hwf+VW9A+Ku/w4LeDOBv00jrDbyKWAAmIZboh3X38tKQ4Jut1fM7x
BPz1ZnN0nx0d7uu3rPzwHI8TZZqQLX1kcoijgmwB3c/2qMxg6yZy9IFJ5GlfoKBAU/V9N5nNWfJg
mq3p+cFdngBTu6mSxc7mHjqvSpByPcTyjBgr/VU+LM+MeETtKfZGJTdLfqFzUKno6uJLTgAA3nV6
U0aB705ibuCj6wSyUFYStgQ+pvMxCB/FkoT5/uY1pAVrGrGCFOhJTTqAV3HL8aIyas0G/4gVsDwi
mTMZXdLNPSVJ39nFol8VPj39GB9mSpLUBRpbm0bzSbUcS4xgx6utpoR65RI5OReoJ+QGnX4VdU1/
2fHYpWF0/x+CaPKdCaFadhDgd1WxM5fJ2qt/ZmybO5BF5iUceIiD30VzVwX2ej+x3BV1gDAwlhRo
Ck3o6e1Z8JbXx6RzTfLpDlV3qNAfbQhM54gwIEPMvjFpbAqLYYzPj/k5UhPxCtQZ4SkNUTPS6k7w
nOp/rnuRY+D8Wnw/f7/QF5PoBEZ/vM2QglT4pZLWYE/3GXnj94o8NhZigflW7SdZRjpKZbuRLNE+
mh3NwD+usr6KG7fCno7FNKdSKlEVsbOii0lzfR+mIYC5B54q6wdKpI3dFndasyhHAEl8SxreCe3N
qUqhLD6UHdEP1KrZ92ID7gU7ixk+4hUJc047SqnjlFUvLgYC5XLi9zPblHmBTbeVrduTiQMpwnp7
F3KAEqz/2NkNJ301E8QD6U+9gjjmRDLHjJauiYJK7+dv4tTJ2+ATl3GCRnz1BQFIpuUK6N/3cHV8
kKy69KglM6z9Al6daEOZztzC+rsR/54Qvu8rncpW/unFtzQaW+twMUeN0eoC8m9Leyb8w65KzPew
OX6INtIgEQFc25JnYkMHbGxCArac5TjcfQQI8GJhxp7M0zuocNinZdTgRXc/SgTrKkSdCXiWB7ud
TdfetS5hYVU6/d3snTFb1Y+aYPc7FvOgf0BocVhOSc9co2yUqzQgwny9MMarZSyeznsM/ecRLL1J
K8pSxOcs8Yy3wpjcy3PUTEt3EcEFg3PMCJrfyvLVjyADsZ64xIaLy9gQ6He9S1bgPoVGXDWBIiLz
lVM2jzAsG4oyHZZrUBj2385cqb9NvuUMg4W8BJGczgF5mO1sXRCE8hrKOnc5C+jQOVJL2TWAmd5J
mH4MFeYVNxNO+G6fWFNRz/9QB5dqwzo+KArE92Nye5fGtd3QKSQVWxm/6qrjLTYycGhmMWEsSie8
AgDyW3U8obxoxecAGdtQCskOgUoyH1WZitKAW9QsxhmVI2BNnTJJjGPC5kz5LcEd4bTB7Iu1HYeQ
h7mWL97pmDMMsKAbIzpksVnwslLLa0Eetqwf6sZ+45n7X2qrRmANe4j44CXYZepDwcTM+TUurd9B
AApREDWvmQYAFX06k+jEISv1mKSWmLHTJ9izFNnxVUO4FGi3+pAGL5KqGVSG12PYf5GySphJv/U6
AR7EArsaUnCol0813mmnIB+hUB0AKx3qVQU1Cn5vNSdYrvi97MObI2byNC1+R/U3s34PYtWsl0Vr
hjm3ZM45TiR0SFxBTl3PHxGLGz2m/NM+ZDbZrppANefXnihHkkDlvprwJO5prP0mwCLk441Bk7cO
qarzME5wgVpje23KQ0mOe7uZ520uV2RavkKcOyDS4xBBxR8luygV9+pGBCcoFQ6qmoeYeLZxhCNp
slHo/IntURdZtPT0NAV881TJVQL8usMXCpIgMoLUH6UlQOEk4zBYl2rVftx95JKui2CCyWy22BbF
UEYawONY2QUuFTOa2LW+i6lc3G740DMJRpze5k0CYs8DRFnVFjap6muSOYAunImUZGrZBUlhPOk8
zf2SrZ7ViiU9H28ZEFTiglLh6Ggi35lhSF2ESsl/IYVTncxKrePIkvfLddBEJyyBgZ7vAzNMKTWo
OLsm3rtMjQEQ92ySewwT5FBnf8V+G2Ypn9pybJDi0ckRgzITMZkvLMbcvH5dUpoI3jVmOWaY0eBH
8EPfjeIcJUiCej8NtAoJheVV7mI8J8LedPvHU5e2L4yHbuOGMaHN1r4cassHeM9G99OqfLgs6cVh
DG++4tr+GJfKAd/uFDpNhyZl2gjPuax0laymCRdqaNG2Mt2+hnbB8POgkFPRhUhxWXxCUQjMTL9Q
RLylCsKu51lAJYwkeMFTdTaQp/EGyha1dLqALfHPflLHbcWY0cQ/05k68RvRhgzTKnhBn3a8uAkH
8HhsJDyo29deF6HqV/Wa7i9yKz6LUM+zVI2HEu6rtRAs14Ru0Rn12IJJewH0Qs9cXISTA7KVlh8+
Wu3M02+CoKO80MEWwqa6YbeiwJP5uYvqsTImDaDjIj186aS/axCQ2YFrz6IWcfU0Pj/zw4Ahrhmg
miiPzXK0cbxaStwhpYhlkhH+5hSLe2QgWxypIIHxVf9K+7EQE3EcuG5IIn174PmahQeZv6WusbnF
6dw+c9uQkI3bivguDL6OfUfROewxkKxZm+XYuLSCSkEPHzuVkDzsPSlQaDyrKwyvqhL5pH/Vf+Pi
3gkkXLW4OApHxyiCt5U5mtHX77fNYRABI257gArK4sNUlNhLOjCm9JiePxrhwsbSDfq5IvJHDEgA
GICI+eusdQ7GYmZUvbG0MfGFKoprhOy5tvk1eWXGSfU8GGNgvOgso1JRSDx5Ks4A/uGUy/Mv9JPk
HUdvVJiU3L98sItD+WnKDGHns4Wr1QU40yGetj8XefCgHllDkQPga1PP3cfwUttxBMyMd1X8y+P9
Et+ulsJ12XiN8LHZEtLuxbgLhGWoh95Bm47xR7Lgd3M3kBFZVuMwo2wB54sxYTLc9qw1cpyUXmKd
EaBExQfBJbNnM5/bU/8oaOtulkMRFq0x85sEW21+KTwJr9SUANQ0s0GevwpyZGLxBJ/1FUsbR0/O
aX+fjLAAHNjZzLRS3Xdw1MDANi8BdEOHxXUZN7dDt4eD6EhQxZz5esnqWLxsc1bZhrC3AAoedVWM
2aNUjSWTd2BsqTWpk67j/njgJIwYthOZc8iHsTC1/9EljMpEf9Te1BhPlROnFWUgXO4BO2rFzCh/
gC+H7CbeX5Y2p5IuwoDl2d7uX3xBStR/GPugNWCnrtufxGUkz7QVaXqzhQufCH5VtJzR6ACSszPa
fnBHlwaWyqKWVZfSoJ+htWPqC1Jk5ah9jxuhhAAz70J7kJnWeLbSfJe+2GlIuYmsj3iM0YuahNY7
CVvKUtk7eKC4ToJ1fEqsNhjjeaf9PvOju75c7ZOwz2U2wVpAc/L3ItJS/zAW/WXhCPw5EAAooVtZ
hbdN1gjiaJKlqpmOcm8imc5QtWf8g+RDOKU+T0xCJBjsgh8Y45iBfeLDhnJvg9Z657hEzzVkvSRW
pwniLxUuhvlbXNJS9iPlw2iiY8ZSDc+Pm6Ee8GCSbH27FJfl5H7FKvhXIyCL5aMzLNFBOWwRUnVz
il7wqMJhQFb9LOI3cYDxG8LImvJ5SNtGOBNRQAIUp5eWpq9kRQiU7q6mFLKlbU2Ii2ggTUAkLidP
OdiYx6usEcG1UBr8N3+MyA4kzva2gCqfxQ6dU+QmKSfBMRWHoGhNVIwyyzUwVy1gw9m0XDUzw3EA
4dxqr94z3Zv/Qb4wED2piCCAMgQV7/ZMMmyjXwT+75LFxFQNpJMz3OSoqbnPcJQxaryMc6I+NWvP
JEcGhIDIodiswTkgaG0DWRKA2g8JVvHDDPKuAu+L9838oy3UMu0wk7/ZFKH9WKIW0ID5PlvlgWKw
JGHq7Ba/PjT77OWjv1kyuRX5V7t0WnjJIvOWnswTR1sOk0rum1p0jlJqcUYiTkNTsIXX4nq/h2IW
w1CIZBYS6CScHmveIBWCL1/Se6x1HNb2D3AQHCmOShq0TzMDEA50Tn+Yeer4qJ7vpErBa2f7XzMF
B+GPBNBL8LJ1hB2rAYV+oqgkTidNR5dZUDOPwbn4N+ey04O65CssI3Dqk7TD5Ioe5+7D0OGGN1Oc
pNozqxAJ4p4jjdo0GYjCHZtm4dhLrGs+TEQ/FM5pIIHUEvOmGHwiz26MCe0F7k85OuY8zGMH1rTA
jmwnI2CtP8fn3v1/ze2pzORhAbC2mJMWhMnq6anE3A4nQo8bg85vb3cmirqSurDO7KAnMNGsmgqB
L6I3QgE4xgJbr11kcvtUDMkvSaAWUoI3Uxz4WyD/lHbwsQK/FEHqinJZ5H5sAlpQ+GNS19Gd2dLy
RJWNQqY7FyA2Hb/o2hfNqB5OBcL3prjEi5PoLFNA2zaOlT456usp5fNgVKXTkabg9wWTsb3dHkDi
8kJA1Ik8eZx9I2pqsIp5/Jvzbxj+61poaCfSS9qxzE2dycI4MZ89kJmXhfuj8omflEqB6sv91/CQ
3TKWOJGtb2GtlEFTwXVrneONzYYZQINu04mEv2dY71r9vwjfB3GbPlipYCvt0ec2TgAkF/POMOyN
FB74I5mH9jb3ryHc2kHFU89X/QLl/9t0dxqVN9S05SnvgWHCfaZAexmSsbTSC18acHyHL9zMfC/m
YJ5A8QtwsPlws5SobWZh/wODD75RxeytTZUcpewJBTHLUGomUMsWJ44TB8asmCYbGkN8rbWAo/rO
aREjcgoYuXR0cJ0DJy6z9WZLNp5a9qCwjqM+A459Qz/C4RBITilZIdDwhuqJyloR93lk56KJVLhU
4x5qs6LI+MtTjk5sCJWkLKIZwi1eoRCEh0jmtSZ58IKCfCyXT1LnOm+EaiYbsSlfws3YlEXfuyVS
+mtsZDuP/Ea02Kys6k7+36BxP6wxejgWomn2CAiSJ0lAMe2wheM0B+Jold3kUPDiHUjUE5eB2ATx
1ccG9tTgoy00VNPsdTzIZ2B2J15aIBDIASh+PUSRMNV5XF9ckwZu0iiyhBw6N9d2Yzwp3xI9GAcC
MDAZNm2deW0uhA25bYWQsNPRPFxAxUnMyThcu5npdtzAR7DycjChq/qRVmoOy5u8XAnC/ZHc+LpJ
UnaRJ1NhJXmW2JC1r5IfsRSzNgKTNBu/Itpw2zdptHzlbU/y1UmG/rQU6GVCHhBogrnfQJ4t5Q4X
uOVFFISVsXEBbVznDFLTonEyAHaaSsK3BXL1tf38olN0QnuIvnwFWu/cQAba7lv9yogrrHPixrGx
2lOSAEw/QwbdRGWtViOOgDE3BwilokmoPwULRuP4iH3p2E/J96Ps/mUy9Zq9f9vDIfUS8IjsIAhA
1ntsQSJ6e9rmErWCS3MF3ukgEZJL4U8jj06oF/AisugRrFTQhevuY+FS3PPbdM2yiMKQbp0dDQsU
9xHMNJ10SCM8bBPcEO1i4gDmHNOpgfngSvm3WSabpOTJkoD6o8b8bbAcr4KEXVFHAWEXOgjbVvgP
miCLxLOa3Peu39p4QTZvAjeUsEFotTd42Q5xCdE6VJuH/iSvBycmbopFzhWkx7pIwFF63d7Xf3sb
0S7ssWMqIuOPXFQ9FRC9klDgFAnCvH3LrSB7Dpl3guF8Z9j+lMnCyoAF8540z8u3DUIvyKaeTC+y
hbtJn6Xh0oX+jR0WKnCU/NEVuYIWvLZCjs8uyn66VLESdrtIVn47f5UtlMKpnIpvL6jaOgZe0wGF
tQpxbNBFN5TLcLenfVQlAGa0WAWk2ENYzVqIz4UHjtz7iOiUVgzMD65XPeFVdsV0uB2kzfAar0zN
c0YslFScVC1f0vIvoMLzdDL9paGcBZI1buYsOB1Y/lEmL5FgTiEu+wDBdHCJELTcfOeMWY4ex9M4
xgZmzR5rTI8SFh3UZOrKYF9fpcUO4ZfN+36qt2tJdZv1KDAO+1HGmKPjNZuyLLkOdd6N3G0J6wDK
4q1HHiZAHVzG0w7Jjy2u7nTPTkzUBRdvCqzln6aM4obCcn9Pg6ChYC+YT+HcN/OoqmWK93SjoUMl
dwtX++FPzLbmTK8+1qUTPXPTsMXpSALWQeYsLUi/2ijT/Bmwf5MrsYIJvczS4mRGd3DPdbPWse+l
U3TBevF6uDNvv7UEhSVgf6lKTH2NJhxX5+heZnoVQX5lLgeyuri5s90RAcbdz6x5SuBt3eNIwtKu
TA4pBY9wLzgbTnNqGGOvW1PDdmAs90d6PoyNmi/EmSHuKRmVyzoGgYm3UpYIuQ1ZAxgaVHfhi8O+
Yt+8foE8k4frzviBIEvLlBWoqQZfOutOQdy/DboBpcpWdzzuVArWHxAsDE1uxLFYlxUeSWZVzEqL
83wNSBeJyG/RvZhkXDFLehxl0cN5OMz7gY2CowYXNh/nB/DGNXXAWTCGgPGE6lhTP3wd3hLP8dsT
WguFR16137+w6IrpFkjo70tREPne05MpFAWeBf75FnigtnUbVl0PNT08gWTNDbYJKHAz6HJ3CDLa
Cs8kivfL9sbcKwiozpjf/DJ5aC0CycL8XCv1ALgqHml5G8ZxIyjhVBagHh9nSZqhB2WjoKH25NIU
1E7//y9gL1mAk8sOCojtAnISHCjbmts+ZlSGuolT5h996B9oh9bfnSikHbWo+w8UWQayPPyWTPfg
goRgYf+CezvKdOnC2amx0mTAnPEScu5uD03dVwtYcwrFy2AmWLavCy4tKznx3Tim3yKA9ZI+pBZW
vOJjau61GddFvjRvn2caYHTAAj27mLdhyiwXoohefjk9ETHqSavAr8q/cCqbRodhdo9FsUnDHK4b
52Zvi0I81Np8w7Y6YvT6RR3zww7Y2w8b4wkqTqwqMV3hGbk39tq/0yYAniFOuuOiqhPDlN+pWOLc
M8NDj5jJ8/WZdeNEbRuHch3zTGBYqaRTS5Qquwqlps6Q5yxVhM7YoLgumGrwxG2+DNWbnX4HGamH
oGJsDHhUfILuQCr8ZYJsM7Ar7HZUUbw4tY3/HklGuquEbkVNGqaXXM6FZijswlkEl6cAtmDH8ED3
V8cZ5nuoBCMtv2qVu26yFoFs7+RR4Kajshglnnvxbx3VDziWGIHYkvtJ2Zjp120lfQ/RNXp0/XAQ
GxnouZ5jc1xW7qYL4wSwg+HZh+4Bxc/KSXYocGB8sbhIveGpasN/6yUjOh1Aws4YQnT28AflmLfM
NHrnqmGLSEIGZaADC6A7NMy6q9Lei7EIEDzkty0NbpGX6AX3jUzi+X4ZxjvQL99KLFmpooW9cw4j
aEMvuSf7lBytFxx4SIwNMhjV5nQHOtb8rirSHFnK/jBpQ0HXkVcnifxbYi9dWuHk0QklJ0rFuOLI
cmHQjfqDCBFA8SqUzanNHtqJJ5VAIUr4hEomjwsKsmDrMu2qaZjaQ/7wqZh9W/fy1/Gtq2fIzq6s
BbnkuJ2jesdF97COSeQ/geCUJhHi2bZ5PBxATp4TFj/8F1nFcVuIf03wVOBXUN6O8gUbRKI6b7Hi
Bc/IBW36SmhQGYSWIsCXV6ZCvGLpdvRFLqApAcKdiASyXuaxY+aVuZ2QBlyhqMinykVKKp/V0MtX
wffVRQFoVUC+w9xBYPbKVT58VdqA82xqeHUSesavFwxQ5H5kUCLvUzkPGGmxen0QH6QgXVfpWKHy
fZyRT1T13EmSor149aStqJPCjmhDWTuCdPx2lR4qWlkPxGe/ND5AbE7PkWN4Tv8kx/nhb2qbxIjM
SRrObp059KuqPHVICp5KYjnzGlabv0UWh8/mXdxnap1rraFW495FBRNQmIQjxFvmde089aSeU0NL
Gv4TMZ7wJIjFVRgRI2wC08y9SsM7MLdEkndj4vJ3Q3VVabxusv8HPkY74epSDchO7cK0W8PMhMBJ
zv9/BOqPwtISD52mffFerynKpI6wW+nCv96QJetz8g3bADyXIMv1o4lADL1cQotP5+Jw5i9jPqco
XqYtLNqkwQZxBiTvVwYPzDjIh44JrteynAIHBgLgOx86QfTNxpvOo1bMoxRIIMHYEpRbZbqv7pG2
6nyL2lg4yfAzRRfqiQdtmbH+SzsMoqi3q7nDp0SGEgzcsjGBswKxtkkdsybs++IMw6kONMrR7xRB
7Q7Z6bBGY/ASES8d+o+IV185m+Ll8Vf3V1Yogr0NvUZYLJFqAs07kupLbTqr27zw0jVJNrrbxnar
atWsoha/u4Z/aCowXqLwoT/3LzcMbPQQ8BGxnoHxleqLvI94Wu5dGodLfEWzFDNyF2iL8v2NUy/V
Skp9Ka31jTPso1lZap3v5J/cZfzlqBTdAgBna9s1bSHSzzRp++V4lZblNM0/+o8X8v4TMx8t8UqM
GLBZzr5zBBuwNbCZLDAy90DzYaKZ4bd9MvIrQz1WjsaWRWjMWHCtXvwICE2HRtjtiULS6nrrq+Tq
4RGLGL7Cj/6KW3IT0hfPL5zRFXq9+LlNd8Xela0eGPhT/h14291uM+cyaGVbJQvu0AoOXdtYAMQy
CVOBFNBdE1v8CG9oLmW/qbTeyh9YVEOzykY8f0HrVM/B4EY0MXVfsNYviqRciOHa4iA9gDI/Uuc5
u38Xz+LyZQTh2OAl/g+/81DW6pQ1+bZLkbC05ZgOiWB/a4zwje1nyTQeTVQw1013+lrUDo1888oA
0iNkSPMY1QwLpIB1kX/lKzEUnQOtZARD3023e/O9UPgyIKUr9Rx2TmBLLel/JOcBY3ZwGjlt04xM
q8c/D/UzC4pkbKdFIAxanFwOxV4MCnDTinw+dqlrl7ZKI5t9gAmq583Izy+bYTg1rMmy/yBCytk8
scQSOADhhJSciYTQEoqSg81tQki89jrMoYabJuQQx09F99oHuzeRWLLvlq+dyNKm7S4Zv8g4wYJi
epWIQIec1ku8+pxKI9XNUs8SgN8h+NZJYiZeAEDLoVZ0ZvVjBVMYtL13l+bpnjoEXAVCNypQBfXg
XfdPXF7r3gW/75wz2LEACBRmPF4eqkF04YVD9R/6ncjRNO1xYNlPSKhqUeID2PiFPG8s7nkBtDAa
Ta+VZXtRcn8nXRoAtygOszQPdRMWsC17nj7HOCj5fET6hXI1Ujd1w+VpH0K2WeC5vjQh5ZYL3UoF
ODqiOWks8Ccus2e1k2utenoceSP+a72HMDI9vRpYQ8bexxSI4WwHJDoLFQwk4ezmXugjLnHP3tiH
dhqc7pwsKFEFRHMnzY7JCZHbbmwLimSHv/xztcuMlD3viVXGo2bunsiih56y1Jt98pCOdmiFnYED
EGtMScLkPNCl9GItctRsKiRozJjeO8aJr+1PdqsTpxrL7RHbruyrx0VZFd/4rOMVXPfoFpa2XJzA
8avGilQKAMHHb4glp44ZwebIj0jiQNv1kMaIxyNJhFs4FVF2VeKaGSzLirLexHvu2VfC5MnH9eeU
YeCIAmbox5o/Rc346/5ZYW1UAHI+htWME0fYE8Jau4bch3yz07kj21cULJ1JYc+yXdY9bK2DKrAy
2Zd30WYVc/o6hRI6IUazJoRm3trabJHLWgtFgnet3xYv3KTg9y9JEqrMHRdCGI+8vgf9P6XIlTrD
sNanJK+jeXXKTyFxlwZ0IOLTMEUx/gLioWQIePTf7hitPmSlzqZVFgjXHCu+vUEEbAWeOsngxgjm
JBMAwyCpkoH8ElxDBc/rgeqFhNbOjwgCLP8KBrjmsQVIgPYhW5G0WJgBVSUtsn/4LtdDD/nyie8G
QF92SH05nGAUXo2S8eWqxvqcSh7wXSC4zasKLwA2neBGOMHHEM7ogNTJRxHZnGUPpF+dFGvTJmm4
k5iH9j73ck3voRwvTykA/PIHugwHl1EsM2jtwbMCozAG7M4Njh9ISIbhmwQ6Jlfw2TsS906WIVEa
h2u1ezxqblOZ3DR4RAKFabT2J+b8D6fzWbOzgO7lAbfiUxsD0hjU/WQ3iL55CzX0wR5Y/nU6nG5j
mm8t+C4k2UP624yZ2Ov6N8VpOHs/Qk9XcfOjE5U3AUcTTJEgW0bF3NsjwObplvOHfQAz6EgKdXTa
LyfTO/1jn+VY6e+avKpv7Y4nZAIEEC2rK6qu30IsRDyHZc2vaTlBFgn2vhH25QTBQX91jc/eU0ul
NRcszUFtth5NzpPBjNRlYf/ZGnXS0EzdwN4d0YYFL+UHgSZUzTWthX3DnUfgsbEqo0w7FUdxMp9m
7MuuYu2QLuUPXzr/RBpNmoXc0vI1vPc/p2YYw6jrt237lnqJ5bC1FBQFgBQ0VnUgV9t81TXlXeiy
y5fSzoiwuV4JPDBwuKMznNKz1MuwyU3IcO9PCwODYpyFaAtU/oLkBPM9nwXlLkmS47khpu+32/Kw
w6Y/+EUc9vwbawl5Co9t3wMG7UJWUVyBAg3XsYJyqjIXkNdSSgMKk1Xu0ukMdoykiyCcuBfpvLHK
nw0LsD67DOKZoGzw4tUTfMdRTRJ47S4o86jqc4QghPRuJZ1Ws7ZZgJWzHUg79GUiCBAuAhDRUaSy
71yNNX47pyg1qZJwXLNdaKXON975Cqx22PC1yygSc4NkVwx0GkGGWSe0qYyooW0lNOCbPOFTPtZ0
n+sZrOvwbh89jT5yV0w+1VMyl8Qt0rbrfVVFS6dMzrztKmE1+hUq/3sT/6dFlwOo0+9kGKm2YY0Z
WcXw8larLCVGCAp1KSGFutkZMfhP/o9oNZLTxZ3TQAiboK6Pju9a3FDrWp6IffSW3feqXFYtWMn3
4jaNyiExOXTnQlvJWUHhzqgA+SJew4laH6s44xXrtos5Gz+Z9Pmdr9zcAyq4yP+mAM6uxGUBnSMO
ZszGe0WQ4EU7LvUREIzh/yjdy6OH19t5xTqJsVFI7SLRGiS9im71zGsO0Po5PDYUCxBB84aK/ZcL
FvZR0GA51UwT2nSoquF6zM0XBfoYcGPj00ZY7sfYCHQ2EI0K7HoCSFB1E4VSiHJXDodSKnLF3gp2
zIRw7Q9W5blKV4gQZnpXbq3G9WCpGvfXUUSQ91yFrr28Jba+XXRx4DaxPPzeGkwHPSRcWAhe1bj1
Gk5VVPk+JlDw/oZDh2Huj/cZHVaexS7jGTaWOU2/FdUYfoNORbkpQHiLgc0goCGlZSAG+CO1nfSx
fOdcsMM3w1PQysKN/8krXLO2H51LyHpMkyKFafrYDwBHpR7JslNVrIsee/79zpc+YOqWQAroVqpS
lvaCS2FNWNy430V/l2jPCJMGdazYeL0b4Scr/f2NmBH3taRAdyLZVX+6McZplUhNFFuTL9KLvuXO
aC/QaK26JVDDtCiGX7wiEOH5gGa9BEhkZaNNb8gXzpq0imhzBWAV8MDnkZqUVZSmyMWXmDshxgzF
SGHifvl6iSl2E+5WQvTQOI6e0ZDraSbR75AHaYOZI2IARhZzksn/1IXoGdUFvmoYF35r7DWrcpnN
F2v5/4NFHenribjmXPbQAVeUvM8P8CW9lfqTIoDzSTiCwJ+Swobqeh3zT4Vmgo34TgC6yE3xE/jA
ydsnJG+L96H0PilWsN18252XnjxgfXpeCkleaBybDLneYJiJBjwBhR6CO9xViGzFWLSP17ULaJ56
+eW2WeonS2nkbmjhWA8DFWgi2h4ExSoZZy6nZYON6RcwP9WKdM/IbI3PCfBtWlFEKeYgGO3ZSpsm
Ta2EZMDSWhwcHfB/xtzLROSU+jCbGUvhK15Kn3eI8BrMfebz0Ejo6eESomKrsaLAVd3KSV+XOz/G
MEJcRZZOMp58lF0LF0y69UDAxGZcfLsUdFAa8tzHLt16z/23Qs6raABlJbsyYS5ZUY/gtuY2CAmH
tBAkus7vHgkmf8gHSQkrfc/ei+gd8IJd/ctNFR0FyFmgKkjhlghdO0r37CPZgkvjK0lUrhrAFqy5
+ogN48I/x5KAwvxL4e401iDTaMH45ML36Z6wdrGRLTWxDsEEgH1nG4wSBpq2XkGKA95ig+EhY3Br
dbTXFlFPWkpLbuXma1Y/pqdsCIDJWGAMqauCt90BT9EWcGla4EXjdWA3TDZrey58A6j9enjvXH3p
t4MQI4JpvA152S+PNeRomy0vvek54KW/zFaee4eVUSFhdRGnV2OXkDz6kxux1JRiJ4cLc2OZ/wnX
7iTsILDw6Y5BfFOyhAWmJI9Uafi8dLRfbKD97fek8aH+0iuj4tZeVZQY2vBkWmpjdgc0jjy/GreX
INpA4INAqFaH/nAfMSswFYuHxQEPXBE2jV868HtNyouieuqcHgpgpwsRWwblLewgklstdWT0LEeA
xe2vjjS9G2daa0zvPJQcfQBXDIudBN87g49Ph1FwK8RjnbsCbgIXUagh3S138vAWKrS3UfXGuqX1
JX66yvgmylEhyHknwFuaNI5W2JM9vsB8HB4dAWpzxSVkL/dJS9zQe/qkFjLwY5gB3NooPi960PbC
gQvSctepEeHFGVA2bNxgnCACFeGVKKarQTo2MXPMnUoN4SS04rW+3i/jwY4mgKg0Zh4WBM1Zpqnw
bjIomSeARKyz/G6CkOj0oBzEJ/bBW1Q9EfRyk36tGl0Du9jMmHid9nTpkOODdvVtw/O0t+MBMYoC
lfJxL58Azj/C3ryn/4wd6BtGkJT0TQi6AvwJBtgVbkEsaywQEmiLiD2nMCWKuSCrNeoORYJSbzGy
xZ4Cw6LCSn8Ho6bZ3vSTywUCMcDpUnQj4TIWsygSm+cnAsf2VpSs6eEzR+0QP9vq615St0TSxuEy
yyaIvOLlKFqE5zOZ81iYg4SifoUkrNJQwYQP+wts+JbXUyx84X6dYhWokYMS1k7NdqCwZ/S35a8O
sUbqif2L8S/1DYOp15geaYCXbCip4Ncf3fPOy6zKq4/un2rqOAZ1UeI+vruf2js0DuvMIHM2vTSL
CGajPgF6OdsYD5j16+P3qxuY4sjjnCTArmBZuB+E9boQn0yz52Dn0l/fP5dvheApN/uxJhlZ/cz7
SSSg7LkigWWui9dUCvlkTBKoFSh01oqPf7lIGfqTOMc4h/mlhjK2X3x+QHKreAxhPbNQi1u0fq0d
xTvbxh/q46AbfHh8Iq7c8mT59/omOmTEvVD1jyrLdXxfHS7iRMRxz/LVgJ/RSZ5gARrZsOjH9Aa3
7aPvzsDEKciPuc120cPHEy0LLRblaLu+95eQpFeZHODuYEqsf0lMvGz3eV/M8w7on6G09GIfZRzU
n5iXOQEyUFVqYQkRMB33EMxSl/uW0gxnwWLfTqacgr4NVGQYfgiN4PtdaSjcBIMVR6SH4vHWssUd
42frrxzIKn1cygXNsZMl+/Uy/ICy5iQtNteM4YYxYfDb7gmMGMAbGD48pS3rspCpx0hm8R/i4hD1
+kYn9NXkv90xPRe9+XUuTyzWo7yIha9aG9+bNnTZd2EykB5x9EWjTCTDfskNq1WEyZWYzT8lAmgY
gBAaTXGAJjBhp2dMo64YtiKAA7cjMssHId5p3FNfJNaoarN9KNM9YmgOVAujJl/wi71fQfDydr5G
JrNdvCC/JWdM+/8F3ANA8L2OLl+a2A45TrMRD2PD4HdY4OmtcltHt5uNe5YgrI5k+3GtRNF0wdg3
GLRzhHqXvMKy+Px431kwkkMTvqU2W/hXZZRlT272JyVy45QIf+O6XWiBfyyvI7u1ssXIwSG919i7
R6x+Zr1hDIChMagoUnhy4iPGMnYMJ9yl8axybNUvP02Z+uc/WCJ1rtDkOG7sk8QdiUT+q51C9NNK
v/HsRPjNc9/o9EAT9gsKnVyQv8J3mhXsIasUluezK2hFHcUCinOV6MwffaxJJK0avsEz/yexIC/s
gs0Q6xoaLk1wKnTGz7w1/IolbUbk8Ln2Uc/VICwrXqY0d6jMkqupTLLsa7h6K3Y/fgjd5XVHMEzh
Y7FDepJqHDKxG5qIwR119rDOdgMKTSzAnTI/uRxM0MKDWNCvX2h9hwIobAFIfECm7K9RwH3Gtk0F
SaoJrePgD42kiEgweqNqGhNgzm3WFSgIaxhoSeK7C3EsIM39wXLpL4cvC4JfQ3aDPQyYK0ceUkS1
mC+rJp7JSrNsZPB0RU/jT/MiFf5bZw7AKRsIKAzaqqoatgtoPJE+PyfZcqo5FS4TfjDTzrTiO/H3
ubYrqEJY6G8W0KdSMPXwTPGrAl9E0d7d/MAKihSEzatpZYHzKmkOvlP316+bwpOn0nFgM1oHt50/
f3+Lzf62h0ysjan0+V4Njsew5PqE8kSNrTqHaTLVyISIMbkCVVN/On1nM4uitAcZEjh3aR0/wtrH
PLjC8cENwClpX/HjGVkiT9qFcwZ8RRgP8sTXdw8BB4VpryrfmPWaXZyLlZ0Y20eW7Ri7RfS6ez4S
3osn6BzDscRNVLdgK2F6IhYet2r46Q8upBzTR6rPsbvJ+xy6D0qudiI0BrhXZ0GL3VjtYb0VlzJF
S4Q6VObgttG0D8nsspz+5drBgMkOFEe1oreX1K5oKySA2fLELgrxsOeP/MXwKvSQqd16Sb38mf5r
TK4qW3glBssjo7eMGBol+JipratdAH1AFlyOKpuYX33Ry00hpXyItq+9K+hMYuzWX+ge4bZxxRsF
aO+1LblEk76WmrfymKXLxtCwl3jzTkve+ac7zPlpIwcY9e67+8rafExPaqZmOpzRO7jzMU1jJ0a8
RYI0BbEbiWx8uSomAG1UMlVvROW5hJ9haHmDzv/WpLfgGDkGBFrOZmquEwIVJrH4kOh5T42KsaCK
/Jgv4kDo93t+VLuVX3B48WV/5FZgC1wavWiCa6TNpp4dAlIlTmIydanmOCdlW8nFYoHyzyPfU5In
+wLGiTct/7uRamLUtLtZbU6f7m0WxiZVLC1mDFCTXNbtSg0x+HyFR+kzTx52JIcjYM4ER5cHqO/w
iNneGV4Fzonvbcrs5t0nJ5W3MzGAMMhKz8wCvp6fJcoNvTApOLGE08NFkECwYulCdjCqmCLI1nw/
A5q3TN2EL22A+FjIvd3pQrt9uQVBultxkkbSxGDAZJy2BgXK2tAsDj1feT2xtF1aKnWAPvIHlOin
AbzDkQ8lvTlvXxMPOXUhUO/lBDxkMP+Ko3E5UV8mPte4N3hEGmNHpwKNY9s0JPeHiHoZRA7Co5A3
1fSUTBFO/utK/kTJR765ZFTlbGmOUNg9HnlGatGfr+SbjgSwoLVk9M/kmOu8lu3w+SVhhDTMONA2
NmddRAYIY9jCtXZImdOctvk2qS2HfU7A2mzEl76F6GdpoFtyDtG2mUDC796ISjAYiOGpC4Iw1/5U
AHrekUpbltkZ/oO9GD7Z0SREFcluh8gX5KVo1113jL/gzKpBQlGThhAKZOIEsmup+zCZyjTimycv
8skOVnZ0JBW143MocFmIFdBFI7GEA4FJeGjoJeOfbihMLs8d/uiaRPMMJKIzXoenti7tMB9FZ5QI
Sx/kj9Mg2mgYU52XjsJg8jQ8J4SgOQ4W+NaXIogwNOzYXYi7OIrJwBGkTE6cP7oj94WKv+XFg9hV
xWSn+Qw7uGqgN5aBsc2vD80mXfY2Lo0sAodOXkfPggxyYIHLo40vwjfMBPzmZdM8zSCk4Nu+KDmu
77Njj2Pz9ZTXwb6DIJ7598T4ekE4oMjbJjC8myOs3+j/47F/5YiqYfv8Xq+o6I7SBmfQkBSuf3EH
0FUFtOZrk8Tip0rXV61Cm44BpkarXvr3GVYVZbFVYXpYhJsVOhn/U2ZDKr7qrbaGKbToSp2j5UPk
9jJ66/+ktqfzMtbJZzXZCys/xLCpObchi9KvEqE+BtRw/DhEDUVh1ikhtbh9fHKJPlMLzUIneaEz
+WbAN3olJbGVTSEo0fm9+z2t2vu/rI6l7kjNMOQWsRHIAcQNlDDtsuLl3N+WVzgnxI+A4mSKzoHZ
rT3h5kn1OjuQ7+aCAay5gL53HukDZdj+jfEUZvzzmFDjede0S0OnGhWewcpB2kV02bIvjGzbPBHi
Gr3cogorekBMzhaVzo+bQFXeeOkkd1TDgEV9d35E8l+IeeJpXHQyDwDOlOOmNNmcQvdQX9K4jOxO
Ppg0hC/mlbdWS/DamwnkWB4rDln4OwaJ6Z3Xb1QSfRuJpqUONE1dtTKz88ffg95hW5Ln4owdkooj
j1NDJHDqdD+bNWNoEwnySSi9pPz2sVTLYHa4Ebzu4DQI+2ork4TJC1n+fduzAhY1Oas7Xl6AFi5V
bCV7Dsp2dIoe00CV9Le+jYXK/QyoByz1zIqC+yPvHRoz58ZmO7PqgfZh+imhYDqxbVrYjPBZSsh/
clHMRtLbzz75Bbva5lE5NCo0NOVHWoD7FaqIE6Z1by+Pnm+VI4FMAz5tp33m1QNa7pEdr4mJVkP3
imEYOTMKcNlSUIgd3IjhOkqbie6vp8fW8UaHvYDHOnCWfKCD5skCUbHvH0wV1/9gCCqBQkQkfyP+
EpFx0FfCfxMrO2b9OnL+kWZ7IPbx6SvUAAYmjyylwcPqM67YYt/pHAkxdCDBeJNEtHmI/TXIfmnD
Ngalr1QwPUsB9qW4t9ccDxrM3XrDVe5t5X+bb0xz6DhvayISNZpYEcxwt4TaAMZCHUP5Lh/90Fze
2RfTUPJ02a0zkBacaU2QmN1PT81W2hwYD+LCBsNJ/iVwvv6H1NWIUkaJ/lGJxUEnnRy7cuWJ+3mS
Qpi2aJIBnlKf6C/xjiU2M7xxHVuYiKf7XhNWmkM3gNB5ZYP9nF/ASrwHxj9qzruyCso/VOVtFJ+b
8bTHGS9HtRpTH/+SCtMS/nMcWjIKRZUhGOOcHHLrt4yaNilpWZC1HtoGE6CUavrJTMKQL0oeJfl7
ZyhAO5/F65oBvigiAysKCT6jwRyQeqtERLJWjYib0WABWinsjHCDNhZlGLJ+xoaZxkihInheoC0c
KxOouSmp5HcaJV8b/MXpYb1lSmGuNcsP5viTmWVBIVrUOmNLRvdZe315PUxjQNs/lB5wv6iJtrKX
gzgP+5R/vQYcCnW3yqTos+iRq1CD8arGfuwaOUUWiwfN02mCEvH0DcRxIXWcPgnchzLDiLcdvC31
mMYAxypQwTHSFSfswU3TBn7lOaQ15aNPEi6wVkwH7bU8XONxi0BwV+aX7vJO4QI0e0LlUaCrqoQd
MMmDHzTQT/ne5N0yYpI+ngjTGf7Lu5vLXJlYYbp5r7GmzJFHAo5K4OVojI0dbjMk87/QH0QwcVM/
V2mcxbLFMSWjdUcc62WRw6Z6OTsWaEodNqUQYSRvOhM3DfM8GAMW+kvVFwnLeid48MZyx3a8mD4j
EMBZgabFl7esKys+lGAZs5lIZYnxD3gNmC6aMI1zsGvTDktbva4KlXkxBHAb9m2OQsIFyy/4v/bi
AGvjebkr3r3GZ+K28b8L1h38GJccTIg5K8IfxIeFlxCBXnpzRqIsDreCva8EHaaYFzEGDEVacOZC
jzcpRFge0wpGme469GG3B9FNaJ0TGd5Ja2L8ybucsk2NUvZh07ue1qmMjOVAb0q5bx6BVjqxKJN9
ELYkYKLmdyv29uPI6FbEFaM6Jim/4BqwNeOevTBYiPLF/4GExrco20mWzTPc8jHecW1sD2e/kmlV
eTK5P7gOLwlrMIwpbZCGcA7gF1IThfvCI8OeZPsW2R2XX7gA5xIsoVwT2ViDMqvWrHICKQmDVWfV
EbValwKK0pqzthp3IOwiPyh2xZ3tRx5n/yB+d72Mz1CYGlfQgYOihlu+Owd9EGtWfyaHHmwZHdYn
p3mXtK5D62+rkJ5b+ueyzs6oOKZVm5ZuTB2TjM4CqsYPAlj9eA6I3LS6jRRjcHNIaUzniiy3kiRr
GN/z6aPzjHICWXZD1buiKa6GzP1gNjOcgn8ca/8586FDa2wkqLPGIvoqLM2dSHYDjVfBEZ/Tagf2
IgXC/qIFjx0u7EQuiC1Ge0i0pUkRXpo1cxCSYILK1gfVDNJyi8IRZl2l/RU/fkhuhLJXvjJ+1bNr
/Qsybnbbknw9RIG906iVmgox9qjhagmaCqWU7bOMGyciA1Lm+jqqJ7oqBp5rejdZRHaiob/E4J7C
BzvR42FqeUp4wLRfCyJXwDo19jr+Jm2M+kwgzkfP7zBFeWbNyjMIfbiYQxbr9Bvlh2ldJVMJQl+c
E0/YGqeEhshyoZFsrC3lxK0Wm7nN4HyM+upJDJHDVMrSWmEo1K98ZueT4BSgC+AB2t9kXxA+NN+A
By6Hi/DL43yVnn5RgS+JnkFZ63mEHJMhvzfr6YBIpq10ZvL7jsA/PdKHdq3+TKNhYlj4/2aaOnwL
uq+AtNb9EgJwA7qJOibUQsPplt9K79UgWh0El9venqDxrUNP9tMLESjDM4Dy2QnHkaxf/URxLWPR
5/KQmVUR0IuOV9u6HQtr4Ht3GR7cIu9doLqu/pBk7aSgvynORm0W3NQIv7u60rdvS/bVLRjzK4nu
Ui6E4vnkCOwbl6ryRY7rfpaqV0AyD4Na6JNAQfX4IGAfZVNI9O1hvpyX5I+vjS+AuWPkOHYy5TIg
5lYJhZykrFtpFJ7zMBHgIN7EOtEIL+67VH3uq/LJzUsHtn00yvg/6n3Qd1XK+V9vf9x4bbnJDntM
wTFbl4fDIS7qVYh49CFU2k0hBasxQvWcUgNwTp9XnCkJj1Fz2KdvFiJQVX9CezyZ/ntjQQAWLWp7
baWGenTLM9P/ouMz/vxihbqs8CbpAgQEO0yYpVFUOeUzqMlkeRS8sJGc7ozfPzBR4JyOG/ymFFl+
+j8LWOM6KMdOOkQbHD4jo6qBgeDZjSgm3LIjsL/m5Jj+kq0bodqtFjhfo/bLRn8ommg/Hu4aRuyR
R9GS/V2+pa6WUDpuS8vvumZlMBjV2CMIXfswXBS4RCSm49MRjHDWKgnbgsDWjF80p16gPVfjUSpV
oTWhKvRluDj29mlIq6c4rxAtGngC8xrdAlpxU1HuYA3O5CHsR5tndIWvivcfmYbJE/vY4IgY8Iat
un9Gz1KnrKVi0GsGqMPx4sQOvtL8VuVmY3xwEgkcKOAoBUZbX0lrMMyuWt800fPeBNuSuyy4VJJN
Mc2oJaaNdh7ZUaP18qa0eHdruRzR5Wydx1OJld5oq+eIQ1nsRrCPkxFnnoN40/YE+cXso94AcRyG
5Q3x2YENK8k25Wbx8vfoGGDqyjcwyznZT0vQgThIfFBSOLozHaAAvzI+vuD+lEEcyW9NBbSI7woj
zlKK3cLkNhju5RTQgY4ojjeBxJ8Ce+BjnYBG08n3ljBASbzXx+eUuD8dC2cwhBmmjQ+BQy1QwmW1
08v2WwSZH8K8HsrGyqj5WjubiePNfufmE6X2WScC94CvMkYp5gbESuIlX41VsYnTci5Qq33cP0qN
WcSroU6/jHwWAxnjnG4S963LsLgZDt/k+9EYYpd69wuQgnM45w0SRhJz1Dl6iY2r7m5aHTMZta2I
XFK5k9or8yv/oT/ePaeDsaO34XNBPjsUUN+WtaqGLr2ez3QY8yvP1PC87g2Fv5xRbaqqM50DvSqs
HGiEEFaWUzBbTKtM7JM6wssUjoAZmRxM22lgEQHDSaAJwO9I3XJnLrunyUo9fj6TQR2NEijNKL6w
uaHSNsxgm9wn+TVvOmBaZ/b+bjYZ2TiRVd7QObyaEvRB6YOaph9gBByFjFTGiWoN8eshlhY75KRz
eCvLhm6hmYcM+7xiZ8lBKmX2iCKBfWOqpCAAJp9Mha7oAstGPww6r4IvIq1A2y4j55szK085GpAw
osBV5JrhLqgCXWB6hrW4M/tCK9U0FMUd/AG4uDLZkA4V9eX4caPIsyZb29NjeE82n7xWogOJp3nD
eMzPI4ZTyjVHl5NG/I2+WE4WL1aBmIJwzKXE/+1JJ6nygcEKNzx//ECXove0MQrpsRPlb+kLKMf/
xsZFq0udSdMvBlnFN80u40n2kNcXMr2j8wUpwrZArmI4+NxKvDmQDy0w0vE7eL/cTBCmmjG1kwWE
I6+Faw9kmnh4MEi+jXxYsogpd6ovGo5WNKxCe/IxW2bfaBBFP7NGjY3ZkoVjy2NYDsxZeRlHFzF6
USwuGjiskgiY3SIsjaNK7rvnAodqYcdoqRKg4p7LamHsCGV9ap8E639D22QEi7wNn2dXO0kYBu9Y
mHT4ZwwhLta+FiUi+R6nz4IUndYbmotfrMuDhvFsJ1m9dFha8GOCuUMZ3kUHfe2EQ6yacx10drVs
lhgSOdJ7DYJpfTipVvtJHbseI/PO8fYuy1Qk9hoGQQNVEZlMYooBnrGlq7DKSgzLKFgWXoOA/G5z
KU4zp0dX1oONvNVhVQdSy8U1JlrojiIyeaQgSW0JauP1afvIg7nIOWf6AQRg5/Z2K3NwS9JAODKM
jZutLIayZMdoN1t/uK0Ek1j5HwZZS3hcsJ+gAtOWAD3oEpw/rBMMTL1+ZlQbGoDpeWCzDf855GBW
IrFiBrIOvPtNw0j8pfNc/VyN5U2u66hAmJIESOo/pG/v2/qVcuHcFhFzyaGfxVI1A/Wy6bUka7d7
ipQKp3IFLHLo1BvEUJ6DHirma5kOydF4sCtABAtvjMRvx3zvZq2CGk0sA6GaeMQag5DBh9VgW0T9
X7maN+U/pbRMjqJeUcrOKeZ7yRhtqqfmZgj0MAw4tFhs7QIVN5mUJnoshlwBdKMBBtJ4SX8pDIgy
x4Yu6iPFDm5Mr2y12sMvdpnnvvjSDA8S307ePAIF4QfSY66h4CvmzMZgngtLKoaQFNyAWSXO1yA+
HmHVJ8S5uOcq1Cv2K8uMXWFfRLkKI7TJEbMCBXVDaCfFJdgATHuL693V8SFWcZ9F88u52I+cttAM
exORq6yjbecpnpIu4CY8zo+S17CLUO24Da9su3LmobuTOsDPZwbce9kl4VAKDzjzLhGVU6+k9lla
zMXSTj4FHpmFmtLpVhYKtcztFKlyq7CmjTiNa2JvfmFEAMGzGYvpTV8/iMykKZOq3nIMMIPJbe2E
leoE6owYKmwvtARGtLIp4AV4VXcNaJ8DjaXd1clpRStO7PFlrOPXeU89uuLwuEvEBAPNe6oLOD1R
OCS/LA0vGZ7Q70O2r2Ca3d9Jq9GLiCARLJDutFSM6PGNxyulnzN2OjtWu2crdvSOPuU0Es6f0OmE
Ze/qF8U/LuXy0xOQqYlS99qIVaNxsVcHKBtxHyLf+60uL97ZVHMqkbZ8LOuSgtVluZWytK/fhxd7
HWRw7ifwjyzm8lLtdKudhtU0OU1oCSCeB5QoDF8RDLilrQQdQgiUYCPT/Gf16wtnUQCQ4+oCgH+Z
1Ke0aFgMD2qAisjcCRq3OFEuDpuv4zYNHTL1dNUHyjfo0YwNFH8F3lCMqGYz9xmeAXAVj7hGD4zE
cPWQgimwdteQ/FCi07J7+GuWsbDsuBgpjU4SmeL3lpgN7+nd0Z2TO1wSi11ERx9PdvZnNTqOOwoO
J5tOqFVW1EyP7JbQxcBunkHoWmdjiJoFhADkjb6rghr3Tg8748QP1Rw1Fj/uIoPNmpdYeZl6BY0Z
wpW7Xbxwq6hLPtXqYJo3dgno1+DA2tgfIK3W5kgP6VHgfMo8+78v5cNoj2QJ7XadRqfGHsFW/oH7
ztzSGkBkOifBl18cpn8TQfXUR+fHTTDl2+J8Qsr/GqnfiFWLhH5/CN+7H6b8HpwQPqgNmkz+Kcb5
6DoogkQklqZkE+mDIdCJDzpQr104zRVRt+p0IJ4+hbhbeKNvImj9fU/MKpSAtBSXDuLbsVr22a1U
2iMS9Ll9MPwOp/9cmYIx4PjhPHjsICeE/xmZDN4f10942Mmv5gHbdVGsvm7ye/fag3Vqd3Kev7QI
c2flmZzt1J2Xf14Bx2e+D/+munl+sqtNsWpIeZuB27tn9VZP770inR3VUwR9/4BTzoT1yay3qKh8
so7ey02EAjC6g1fHIN96td7vh56GG2wyjkn1+1hwBd4MZvBdREAeuD3ESmqQ4sn7UtyTWYVIlc+J
lvdB4gJLjGTjzPTd2zx0s8PKXoVk0ZcqQXdz8egvBY/SHk127MS2VzeWMw53nZgzS0rlSL9lGZab
+WFvtxxRGJXzhn5gHJ/+lKT8zVLhWVjbrfrLsACAjGkWppKPZJ5wf++OSIqC6pGn1QZls5VtnjIa
3HIbLZuffZbpEYQ4X2m4ytu+K6G3YBo+Ex6TXx/gbMYAqFbjff0KgtSQoJSRCa5PeG3MF1dxYXxx
WPkYJ1H+7zIDeI6tKOss6ZJtYs124ebUqCpHR6vZ1nHgd7G7OzWRWb6gVpmX/H8a7cOEu0vVpcSg
grvaO8cqCIg1dPQqFt1FGNWJ92qvWxrNC8lZA5DlT/APVLrO5u593ILWJUZiQx4K3mrpX3MuOckg
90IaRLL2WordFRmiaIYuZL5XPd6Q3ozvSn3Ka/zW7gP//EiNqD7WItUjrp6bsGpH47AFmgBYz5Rj
fmVbXDWJLcYCZIsbgAEx1jAS0tBPdyRCzrVmyiYqo/fDf4sFFQYqzjRPeFWKssc1LN7CcOWIe8CH
+ZMZQ6rgABO2IzqfDeQTSPbfqWZFRShOJ5AwssFaE3OCzwkx8H/xLuMAVrb8S5UjK4ls7GPWCbO7
rektffCoVvmvQO5g3DkgFYwkgKrc9SsieAwWD5EXIZVXqCniLW4FFPa4w8Hemvvwogr7qWlbOB+G
S6Ir2F+I8IsbPM862a7Z68IZ9PgOiAW2U9cN1Bvm6iUNhyeDeD/Lqrjr405q1wvh9aSg/Re8GHyp
HGz1k6ZAeO4HXeMH8M3ZRCz/jGY/xGihPzscpA+XarZMv1TiMOkK1BI4heQUvNyIBVdFEmrDp4Yy
G2ec+rdyiOqVxrqMLjPFLdkgnpw7nEUQ1kfPiC9BjxFJ3FIRG6WY+M6/6GJ/NLsc2TbyzgCYh9gq
5EcMMOE9cPB8eTr3gLOGGHV6awLLEfWZyzwlHzn0b5f+/NWZZ4f89STrAjE5uyoRDfVblYzGUPvn
MbfKnMcBvHlInIyhhgLnLUU120m5FukHs6TtXQW6ZIgG2P5fkoFwKeafKh+tSY5hv2O0KiQb96mD
jEJZbBsN9OatzaVYVSyvsOknG+mZ9dPnGBvDFuQa1doR0Ey6ew6BapPM928wA7NMN3IB9jX+sxWu
yUa1lIHYVxTG+p8JM0z9oVwHlgDgAo3oMk41NB8bQTb46gpGNL90Qeiq0x1vzzooEvndl3aKtO1C
MZ4ABJMkazmfkJauy95tpMAWsnCXAyH+ToVQAfwTZNRaBNxU0dq5gwvgLGqttypPefHnw46JgqI4
WC0FcBCZwmVyBM/T5Yanj2q6nNKgJcqtgQEVEGIBDu8RlEf4e8ieSHQcCj7bBgUvJcNtu3S2OY84
j+CpvcXuyRuX8J1WTZW83Zx2ezn44Qt0z2uszvgoFwriPJ+kcHE02ZxzmxcwXOhNkbB0j7yr4YgU
zDuZwpGK4gzvpTTAR9fN+ZFYfh8++3iKKg6+OfTN38uHps5UPIemQaJKZzaB8FCpz3JWHeetxsJv
1PwS4pQBEqcOU0aXP2zZx1btfuxwBnEGoyPy36kXQxnuAPTJic8a0Uti/Y2+msUCxQmdx0JzWLMW
lUoXhuSt5ZgvxRB+XOXmdAt00B5uX2Gc/m+0q3El435L5a1LIxl+uOeyYf5ykZo9K7cEdPANDZ7A
S9JVICjurD7nilx0xIrmScNvKE8vsGT96/nSy8SyyurFfUQUgpY/EKF139cD3nsqVV04aH4yYppr
uruMKJW8ypRu9cj3V95N4Up6D96s0H0lBwOMiryR16QOWftNu/9qne4yiZqxTbQWuJweLJbMBJne
ZEsiqQ/OCqh0WRzrm8O7CX1rmPbILSdMYE0CujNWLgkJt0+iYP8DUCz1UkQWnhrHG0VhTRIDWfv+
WwNF9m1gxR6IyiQainog1RaqaA7VcQjLnTgEIxSlxANGNwEVIe3+FD5goFkLcEp+b+e4tBDMNYUd
G5+EnuuXLMNyOd1t62jp3LObtLqoL2FWxKrh+GY8khJXZWjZq3mv/DkL5HZ89qZ3ad4YsYCHGa/b
C7+NSNY4AQ/76bITIbFhwrIEzNLcCJf7P+XsBbV3aJLX/9iRPrvta6Fhwh9QgOgtHo2FXsOW0xlG
78Z1rvgSkedqfQ5qEI5Pd8Cm23iqtRfA2A+s4C8K2DXwbw49QqkoWhMTHnRevI9LfBCih99/yu/P
v69zECp30O0ocWvSh2/j0RWR0szZGFPEiacsTmX1nCe7n3H8fhdv8qR8yBjnYTO0DMViF3olhY/5
zy/3iffF94QXxJtUmpcEItL49VqQ6lI9xKJknz1ltxCN3R2oYdpCOTGEDZ+Jjt9xV7t8+fPJGZCm
s9OkCrB3trplq9IPk5TPorndQby/XU3GFLdz0JH0hMfY13FnuZ0yViuM6DJZx/jblrnowAga0vcn
K5z3yI4zb+J7P8NS8fysAOoEoTAr3eE7oxAUIkhpBjvg5L3ZBsmsDfA2xjhcPOZilWNVXHlFsAKj
Dn/uHRKFtK4mhauWLZ9amXX4h4PKKKOV8LscLzHRKZl9sJ7uzcklJdy8l9KLfgHIvNirbJbf9t9s
7bhrKfLYI8tEhEBWtTR0XrMzoPHLTFdoyHy9ZaCsT1/pv3er62n3eH5N6eQY+/8+yUigb6/FVbt7
84lv4oueAA1IgixQBt0g/X1f1wpuXfnl0WdsJm0giLMoYadYZAwfxUsoRJ2JgOOioKBRB7xRN4uC
qIWYp/p2g6VHjHl9dpLuzfX13dIU4qsHRQcOw27pUwyi/+6Gl2NpxPu5V1eRUyYcns2xKdg8PLOP
2EiO2fQfrnKiY5qSvVHJTnhLOjW4jpcDBK+Bs3B37/nbFn1v605xdkBQXHSUYkOqJoTZf1RgoUWo
fUawTq5Fnv62XM3vCCrDyf9WnE0pciw9qs7KqtY/4z3nToWvjmDKJysuJ55hpeUd0HnU2i67xiQO
h8RR02z30IInt7l9BOrB3na9ag5pGupbnEKvWpDkegvoVlYoSphY7PmfLe1mG15OuHVQ0zYKOhwW
fGEJ3TWdq/paQmCR/zhARm1DyxupNTAaXxFRwiDwdbUENBJ+kXSjYtUo5VAalyGVXB5Fg3VGqiVw
7SUf6FyxfMTNJba297gLGV88TLnONVjJXlyssOub01CDbQmyNl0/QLpjEgXLPIoLQZQc7Glzt062
TxoU2ZfqXJq8C2MXhyHZzt27aLPvL2oEPhi2U8dz6vydhbUgI0XA9vQmeedffuh3uSD0LUFnDGC6
OlSUALmLm81mE3AOxJ3hk2fEuWzzU13awMrItjetXLA05UVXSUEiINpiiRnEkvv8LCHLcYoifRhp
m/yIdZrO46kTyBGzVy8U8BzdPy81IcF3uaHUNl3ZkQnDO98eLanTxTv/z29jJvQQha9OpNUQ7Oae
g46UlxHn8rF6nlCeCISlOYVfxkoQRhlUP5TXCTkwJT/zvE3036XAfxlC5foBLoGcZCd54eq4yDn3
WLPkH9s7LlsbXywwCbpCOTyPF/5z49sC0+0rX4IpyEWLPWwuQZz088ByjCkV1z5BfevgjR1nrSR7
jZIliOVhwvmoICOYbhG29vVw4MpeLvpa/LrEYCXdKduffMd1g/Sg1pE3okEKOPY4Jf2whu/zgcwa
VmQWoUeGgch0NEoOVFG34z3yCHvfieXUYWFDF0Mrl6k+uzn/rUV/gO158OF6g3MmuKbH2enErWou
1a6mA4Xz4ddUhlsH4g2pkrtPjTYA8m26E8KpRav8km9IWFJJ8eXdT2d6hPeCQwyCGTD3z2a4RUqN
HxFxEmKqmRhsLdDvg8hNbHdfJGC+R72dbxwrbhwuvKl52LbzjsjFcu/wBu0nEPqu9SBGkMGzAclf
63EPpdmmNSTpNl9jOyef6CfP5ZhZSJY8mo6SfM4jhxB2F9ZeTtuasy26hyDKzV+TYMf+EVy4vJkF
zCinfTFiF2JkfcreGtLKEZO9HN/nMKINkIWzQ4o+5E897mqHK+Gsw5wO/F1k2U4aDR558TrRYepY
Y9OGcKTV62V8AlnyE60uVwGUdigr8cpz/6LHwx/SaRm5a7RqYctcVrdQoUw1VQCa1GMpvsGtPgNF
dmoBKmKavYz7eCcPAV+bKZsTX4p05Fjut3B7awi65Z+BED2R0tC3d/7QMsZcI/DJQL79MINajZ4Y
JO2NVN+sRW9XhW/ISak94TyTwPHpktPMxOYWnNG4+KpFWXrswpPnUodJ50aNG0tkg53xr59RKxc1
rckODXhDel5zHZ4GHoMBa9adVPDApfb2HFqTEv5G01OzRnSZQlwmAD+O2z2EhIPGEZIt4RainwOr
1HWiYj302qfYFaDZTaE2sxHEM5NdobMMvMEpJzqwAQGfxr90NmraXADP2lfYm4NVsPKn7ABsipiU
JXGW5vbxSoIjsaeqsdwC2gxpqmOYSSFrgbOEWGodYNS3a+wGr59v8Q4EbuOB5uAesAkJ5lFUjxFc
0RaOfxt6q0qGh3v4xtbqAPJj6bl5ibQ/NAcs+02ShfqqxKokl+BZxj5PjhIMx5W9bniQobcFE51S
xPuBRa1R21PdD1X6iVM+ES2QGAXIrTs6nn0MebVyVp+EpAzGWPVydHz7Df5Q+BsR0lvisvz3SuVa
WHzHuyC7wL7KPE93HXhr84u2YPMNjm6aHK3tTnt2Nm9nO6EINbzmGNK5KEhWn9mdhOWMq11ziGKm
Qac/50OzvhijMfH1CoMutk4FLSG6cV0qLFDJKk+Ybvr4EneF/RqX2Ur/+M3cNIHalpGZSnGsm5wO
TIdbuiOTOYNeaTApQnnzeaWPrKWbUxxPNHBLQcB5z5hhKPAotEzweC5u9eRfgctsEmCZrwFwOwmH
g1NBHo1t4WjHemCZ0+NKsgDJ3Aeb4FjJuv3IHCaECQ5i+Aka8K56gr+UtB9IJNEAUvwX8YrT9i0V
OLAj30W8rX2eSjC4Q0ZIeEqGAMB0GdlymBsOpRhQAweSr86w/E99KumBKhjTvSa/caWRWqZngcR3
M2ZW4bfuLTlUgy+N/QbMwXA6MOczIo0npyAFfb9PkPDRWCLB1tvmlERUgmOrW4NC8pC9YxMCsoOM
azpRrjEGUulT9juIkS8fHCEaoGzvTrcUc6/GRsAKFIdkwURlAVwzkkK+d8fELjV2NbwhCvCAZqK4
/r5lBc23trZr+MJ30LobP4nG+mBsdZtkicSD+mSToCFWqr57pG6su01texAbeOCfLnoXDBb6Wblx
ikrmU4YxxBhi3MMNnanu/yt9CCW//VkwKGtFHac8weJ1tK7oH4rd4NU50eGb0Z5hV0eOp4QYbReW
L6uz1dzEDzrb5D2wknZ4hrTkDf8NIT8MkLgOswfxlNK7ErVDAhBNlCGDdmExUltZXXQzpKhA1vvk
WCwW0WeYV4+ElgKQsWcgIFUFdRe+UpRJXX7FOkXVjkzSlE+yxfUVSlWoc4xvWV/7gqYLGSenQSas
HYAMDHXmuNk84Gto8Lf/N9daoEpLj0XBuTLCesi42GghWRxwj2Wcg3F0JC587YqnyScyUd5xykeR
/IvYrW3bM3sImPxciTHlFF8IgAv6gpjdy8oa8AmNO4zsmvadDSISBYfiARTd7sb06Mvtgui6N8Um
L5M6oyZOmFxWyNz7AOdFHDZkXmF2U0u42VizpaZJElzhNIY58lwFO+oS7y7IcjAYWGKsAyDe6DL/
32Yr74/qLfZh/M/3HF4uPkfIY48ZK2F7ajjxe+hwl8FhKYP6FQk6+OI3NFXqFqDre2BBJ7xpjK9a
bs9Dfd7L7KLKpykN/d19hXwgzGuS+IW8O+MBwkJgzH3TNbglNwO/Ixp0taTfQ0YrDlD4yJSRAxPg
WZjIwNpsqUIRdJPHjtQ20qDfVZjK63ymAnJCDskzq5Z2Bh3/eNpFkAvTn8yjPkfjegSBI0wTZy6/
LMcBJFRIrT7DvMa87Ae2ESj+YU5F5BIZlR5v5PF8P8s6HQ/SQoNQPaAjBrdZYPOdn3TN7BAkO8HE
BVfePo+tZrpQ1cvWIMSioV6MLZIIzVqDLlAlaLOQSbD3tf42Hf4ZDjHbU+OqiNc0O2O+EqOgS1nh
ctJTLUnJYVgo3mYGgWAwkcdKPH3mhIRwrPmpzqxwCyC6OF1koPXFtLJwcAl3XoTAGBsIRZi0TaDd
qkb701ZbH0JOlV/fdU2wMCyD1dm0mzXk9vqpzT5oK+7WQiPlaIi8K7xKUp/xpSOMBZ6G/Ps9UrKV
emkGi7G8XHsurV0yaOBU0IIQlc/d5DOhsktnVe823RM6i4QlBxOO943nY/2Mfo+RoAH83V8qrNi6
YobAYNWg4wFYqOjbEEo6a2Eq5yLcMCV7zGTxnUu5VbOFkUaATcLZQGeUwU2alsXYG3CO1y8CuzeF
I9tGDbczOWFmHjUXkGOyCLVz9v/YfW+BC5xCLPKUCLUKVBpkm9tpoBJquV1iO9YRpPAeYOHRWW8s
Ub7NGl1DgFO34bPly6U14+Hv2xfxyJuxoQ7E5mfWjdDBnKeBDv99cEu3gIiWLqlpyuoUkELJX00E
kfNH4RzOtG7thO9f/m1Pk3NF2pODAt59NvQFV3Be08T1AZsFu8jT+DSCqLjTNLc0ECgFMZITsvPf
87cI0IzD6vIPEEEzpoRY3uNVoY1aYg1slQx13BUEFuFuvpVDskAmA6KBlJM7PojCswYKX43x0r5Y
qDZsZJxjTB5CXvRUIT1pYSc5d0ebAgIW3Wgr8jEXbehFs5N+Mbtl/JD5r6RM1LyH52swRrjmjRP6
tNdXTOVAkO5lTdHHVGsDCO47YCH9g5o8cyH+oTAKOPmPfAkLu54brkYQMhZpZ8OuCf/LQp0HTb6M
FDFMIqvVURp00TRfqPv7pnCBjg8t6f07ZRaXo0tcgmsT/3afHE7wtMtQNKXfA9vw7A68H5MZza1w
E948rdpVx+hCxg8NEuLiz9qLAyhpjtGoRwOouvbviN/19NA9sguI9R/QMgaZBFXLQWQ+IcjSYDhU
hCif8e8kXmSYKuCrDKrR06cvv8UX3KNWBTzzjwimX3hqEqnHltyJVazGAmVpNKMKXaSuETWic2k8
qs2r3Xi74F9JkOeGS7yNpFIoKyBCfxScr1WOg4kUhGrT8YpjQx9cWgLX0sdSnYE/ndVgaJCTKXUZ
TVABItYMAlxl2Nech5CNVrwsCJ2vvmOsbJ/CuOFwUNYadL0tDBhQaGmrFENnW8N0BSkuN5WbqFpc
n1iEKdIeVUrjqyYGZ5DYeeSQc5mbbTnqoKEgNQTG22h3p/3B8zPoii0To24E02I+zi5Jie5tUOHK
H8z2VW9dKyOH8TVYaR1Yh6rQZRztcOCFG9xtrD4ClaOYFkfFcf7fFaR/2GEUb9FHvtkAJsbSTruv
GWJKnT8N22iw7Vvo0Vec/R5c2ew4kTIzORmTZRLfu8vB5pSechbgk+FWJLrNzBROj7r/dQuwOmeS
+znAd+0/v0swmSzofxb6O0nE+iM22HjvZK40NJrf1U5E+CenMCUtt6gCG/DshsyYEDrWMr7dnFuF
Rhv9iS7vbsVR/2yTs4p9go4s/ymVo0j/rLoweyAoGmxtl8DbJu6q0Q/Rm+jhFUKz12IMnbpETWwo
y3fyvPCGrPlp43n5N57of/8pf2myuQomhHgqBCMuqvJxyqTkE+EICnV1u5bje4A4sIcd5NtSnGgn
rST/Jgvrlju3wzsOWHqMDdqcayUnpGdzy3vHVu6LaQrt4Zc+Su3p4K5hTWg+rIs6IHyU9tR00/j1
bc82Ql7k81ziy/JVi6mcNkXoPUCp9uSYHwm0fFpPE/jgmcu5m9kPIKfd513eLYY7yOItbfXx31lp
xyyK9+kSgJz1TeMealtV3tst3mcpcy/OvfE7QZ7kjgf/oDX32gcA1TlfSh/35Uzlc2yOdS0uUGTg
qs9dz02jSHYb1TJQOTvBnNhASDKIDauT9etMiVzFaw/yxYeoZg+5f4TNb6E2ZmcOS1bdeS8bDn4p
LGDQTKsPLtEzeFfF8WhjWhbjj6M8C6QJCeCworhuzmyOfHqL85i6sWxW0s7CsJ4WuGOTHN9cEBsu
2Ll0B8w1c1VRWbgS/O9ktGpZiram19owqO0iGvjOGzaE4n/rCloxlsr2SRYAK66YcqVHylnQ3I4B
/8O5mQlkjXpFDFdzPJggtdDWlpNhra6rYOB91YOXxcg7kFkbXve5JOK+ARppaxwF3CPXPiXjU9Da
upj2oxu0a8kM0du119dNXvWNw0gGBNi/j0jIKgfwRGteUwcV2SMLV4UY527FYIHEVG7ebBW0ZhXs
Dtg409boWtvq1CSGAfH2OYddf7TUKEp1RjlGAlXcMGysW/Er6Qey6GAGnfuGJ7a6OIJ/a4m91ZB3
264NuGVUxv5vIwc9Xsh3A15wNI1/TOwxcm6yBeKckuYsSzSwP9aLEyHu7rCMCeCqVKluZnIabvz2
E4Rqxf97KlsecFd4ER0SKj7hapulPZ0I2aW06c1p+aIavJGBDJswCOhgzbOOexi0XWJnzV+Xa+Fq
uVc8mFToGfFTKXwUN5wCOpBwobBPJn3U1MtVqNUIEOvHQve/iogh/FZSeA8pYWR5wC8ViGOP6MnI
q8GD8HbGeXP/jks88jkC12M2mKS+AseufldXOU6r0Owf4kKktgvmMf2HomFX+q2Qcir99r/CGriV
XGDOXSiIONhd/bTkI37VmLRKcScPdYb7O3MM5LwMs3KfdPY9qJwuoWATOO+V1CEjmyuV51uxxCDv
vD6h3XxS+/0HztNCsRzPxQmoo2nYX3moGanq5bChxhqhzZEYBF5laLtinaXpmKCF/BOo4dhT6v+W
jrE9H0TEf2CdI+gfOL4yax7IL8CCuvpITPVHCPy/MBQmXRCLjRAcRIowP+SQzmA8Gz0NAw+M2kub
LODysex35j9whMKNz/pzPNIZp/m1w/M7rQD/GfBSTzLc1wsiqk6xHAX5orPVIggM1EgZ7+l7gVab
C5j7kqix43GmV2P1gqpFdjVzitAueY0/4E40f9cDB30aEMGmThYUCigZm7TGL6/Zhhiu6kTEt8y9
638syqDIOkC5LfZ4lgFZOxwUl6t9+mXcUEov5zkdO6WYLCeqjWFQdvY9ekBvt3//2WcBWGlxGADV
wnBA0os5xm8ekxs9TG6nZG8o3mKUO5QmHoltlNeRx4wFeQaKPU60qdWC639hbRY1flaC1/PZZCpM
8tz2LTwZ/vqfWZDsRmXwcY1qETI1gWC951wNQ33EqnrTwZfVhVgPo3Up6BZgxfuyY0cpJGeX37cK
lT8Adcaps4YSnrALZWxeeQkPSDc9R73CkvSSXdcXuAnumF8Bhso6k8Uel0adsDYScG4SIOyKhGJg
NXoBIfI6GECGCvdv9rBdDus6FO9mv/hhfqN/p/iRs8QfJEoz1DAWMzqkSenAqxPHoqebTamDzSVI
fq8lf4TYZn9Gh+NspAyniVuDZClAJBKN8575pTF1ri6cdxgzBzJjTQxchEYTKNe20RuqzxMFb+8S
tO9oOUUtpnBNtPGOy8GyIfju9wrAgnIRRZfTLUZPQjIoC7Bs+VaUnTlzRrgDXA1BZR09qc2g+gjs
8sWST2YRGE9941g20DYvxSx5UIomuKVE14ntrK7LO1/+ajnvx46KoDXHw4aDRKoBSWLNrze//DmU
Y39RdwFqMRyw8SExg2iyT0r4kpIlOqHfa24CX5+ZHOA2SgdAEqj7p2qX5oTL93H9IEGNPdFZxwsU
h8Z03uYlHtySRwcoZvp6yVHRTJo/gwABSEVIxFxExZKV7SXC7ml7lAPvh6Sy6Wg/HZVbMTrNgiKp
OhtFM2FfkziKcASkeUK66Otk2GxpAmYryXEuU10jRxDi5fzws8aOwY6KyA3uKckZJMV+f4ddMH6F
hYze7p2gH8vy2/uw8MERaxXrnBqoNHUlqZXUCEQDVTIriEUOsB0BuivKXToCbkZ1E9h+X6H9yLtc
tXVmRMRjF09yBPt3Yx5940ZRHYY2Xvo9kip6FGy7ZfBiF5mabPtjQyKnV0J2fyFHB54jTq/LC6tB
vXWT7h8Cd9bg10+tAGXFidQtRPAFnhGOrXKn2VpjFxfMLLFPM8+aNIXh5EA3dRDaSW1mImaIEGC3
8oZLDzEUfFXUIk2S0SlRISLXNMzL2k1uzqijfr21uHa/X1kwau8Vc2b56otwErF+72JLwrvrn45I
bJaoxgRc8Rl2NuVILvOEFEUthPHZvhjpcb6uqADa4y6eOT5RqXpJSpJtpmXESp6zD0BNVl9WEouJ
NZgOKTnW3NVggXTEYp/7J8jyGb+YiWaA+cyRZ4kE0CtGDQlTfd+vcHz3BC5utjIZBLLNaNgkZ3LB
odXdpO1hcCK8V1ewYi39746hhaa/chDsO/35S01cLdRMWncnQNoZ2AnY6KphC2ukBUUWu8SBx+0c
gyktGJI/A8yHujzylcYR7/A8saaXo/JVWWe7T8yXK/9shBgcyMOxgyI5RittbtLjbHY8pXC940+N
fEpIIFNh2JVrZmK9MHLarN1SaxhJcfD5zDhmEREntd/szKiDcPxkE0+QMxhiw2CRpXxAlEJ1E3c0
sgwZye3R9V8EiAQkfTzN8dzuW0NuT7nrn9HwXPXV5tdAh63P/2e+UllAb83LLtZ7+Es21N5nlRCB
8H6iSkowTuYW5UoyD/y0sLUlSPs0Qn822fA17V+WNhzxnMCE0LJ/Kwt03DTWZyx4oTIntO5CQJE1
TdppCeL6FJhG5qz0jTNCV/I16b1CJCrr3qFt2Q0gzBORxAH8emjVxPfrN68zRiBGe5Coew3T1i0c
BhwAC//XiEqdVBMSj8jZ7LWeZGPDHyFMipQNU3CshOxoxFVyfykz8E02DTn8XWb+W7iWPpfkuG9X
7McSQnAios+iM4N9D5zrLkHZpibhmJlhzcGtu9SiJh0cXyQnKHe1Y09mWX17jj4OBqC4jB3GOhGa
4FzFAyztHXpKOBIdfnYR6Kmn4rVg8B47Eu0LsIYKsyQM/B4Y84Gr6DUk4P+MEHcuF+T/UUBO8D4t
JM9j9DjTjM3r0sEvmM/LIyOMGh2TgyKrtcZ8ezALcviPc0PB2C6VxF3PGfnYCKJgIrQ2kJywbRfS
J/acK575gkDazxbIWmcQr+H/YlK6vHqu5/2j0uPS1EdyivgjezmO/MDMwPfTdfAN7foI0e7W75d3
KvTQgQ1Zv6V3v/cUgEkvYNKzPsx2rq4Y1kVB7rShaqWonYVH4Ezlgd0mI9hniv3oVsNjiBw3SqpT
KnUxYa7kJYaCvUWSB39tfaVvle0PxDIc3NUFlGVbL504uAIZPFgCRupUJHEZL9ugogiHa+pCjIVC
DUGNBgk48P+pupQ7foNrLa4wb1OpXAJwg7S8F6/w9kdVWAtZgdvp6SEcxx7R+QlROzINSWPCxFZu
Uvks8IHX9P7HRFp8RodAeM06G5m0hY0l4DO3zp3ZR9woB4Nj83nWRF3VhAg+C0xBFgpmLvA6ejP3
XC4Arl6uW3M06bGJKpnA3p06DY/UtFnMxCxLRhNsDgmcBvvGmHxibVPnfGijhLmeWkuOegHkCfee
Jq/8s8M7vTZKLeUnhrD2QV314l5cI9wO/RsKWUEWwK0bJaH0Awg4QMdSKbQvRdqU7GHJrlD1Qqq4
zNJNa25VZmB/TMGMuGxo27cHbUFt0pV5zBNLxcptzkFqoskGeGX40zBNaNkGPqXncJqRA9jG4u3R
eFSICKxF661w66tF/q6iLLpMEDdr3fz/Ce4wPMS5kTsv3oiiALfPDxgw1HI6tmdld7jvcrTgeN7R
0kkNxX4cwSNw/JszxMP1AWfm9rEkT1CZjwGI1VKZiO+mBZsTEWpqjcSlMoIpxQVTbn/WDikTwwWm
E8bMId92FYPHbbj6FEno/UV9vgR2XLxkSUGAVzpK5MxQLU6yFtGe/Rz2Us2t3zRei12tNBJGCGvU
srqu4Wzv5pPEa9kkU09Pd0i0nyFYRWuWOFx3GpF7vb2wm/vnXB6/LzGl2h4Mox9//0QNbIxzk5So
PkDUmYcTg68LAMX3yN4Oc6d2AtDQvHY7hVNkEGMEecvkLsEYnuG3Q1xFb30JH2t7kg0XIPzeFpf1
NEvNm0JZC+swfWycrgA5rZUaL/JW56bcnVResyIy0IDzBhc5uH2JVe4B7zsOnEIPPh3fqSCFAq9Y
GiFpK2MB8wJDj2+DCA8uz3nscG1B2VZnoNNVBJkkYJ1yah5H2J2sVK2ZqptzdKdGRdJnRI0TuFtg
dzUAtWjUGGGzObCnnCKzGvobuIphIYPaNAYtfZ0/SDzdGew6zr4/lJ2hItySIdVqNUVNsSCzkLuB
FQbckOOK7+IdFw6/wxPG+/REaiY7b8rUlzLEK+iQ2LCrca52+JUvnLPuS7F2yNvdjFaXiqrd2hLG
svSQGTfvmTkDEebC6+bYcJe9Ir0eqe/khO/1uWgwjKRadiiSDtG5sVTkox3EH4tavpX+5lbBo/xZ
vqvGK+KRbE8WxbobdKiwl2YqjWFIn/+mZhiW0urpH8sRG0HQvZulXYtGuxfMXRHUW707zA9E5jp3
4/wPs8KSFjqH+c9HvBQcHADYbR5oGJDVnzCGvLnEhcFxGj6Cd5+i4fYzKJawIrGlohRme6JkBzuV
IZ6vj+0G30IGBpgwjnhNmcJOdC9uegzsd6rUgrcF89jj3QnQe3mgmPNWzMTsV6OqX5mHrIjNpTUX
bR73wLcMPPoHXXo175dzoeMHDUU+aN88ivy9IBD3NOkmBDltuve2+5Fp8eQRBRYkJdl6wAsjx6Nk
qDlrJELXxwrTt9yoMTQfsTVtyjO/l/+s8Y876GmM7GCO9kz3Lnm2eABaXyIbN7hYPX1KE6lyeusy
+M+7P3uMwkTyNe8v2Xj8s7Gb3e5gJlEN96Dfkt9O4TiUuWdX2N7xjw4lZZuppI3WYg0kq/1F5mys
bXVa8zEMIeKNwu1NIuM+jVoo2hic3ILayaNabKN+9E95i0u4GToTf47ykya3LGn9+nZ7M7tJEz4a
ZOG3TYQrL4WtABv1dzJ7M5is90goWavHjhYARTAs4lvpsPZLFVcQrTLbbB/9Uzt6cr+KI7C40C/H
Xnx4Hf+eZRf5BlXWcTo/MAxFJj1We/4QXOTfJtyy5/VPQpJirVQfS1OXTg42yzIUCmsejkz3ml8V
hE7kp1b8CRKKGbZqUftkepwHEuRJn5nE1Lc69q97wasI87SOja7lB5/8NJRTrILFJrVVovsPX/JR
ZCoQp13zBwRYBfYhE8pyYjdMh/aLoxyso0y3TGyub2h0U2oUMGbVCuZSAk5VTM4Y7b+bgrUK70Q5
c6KxjAmeo5nhG+XYzkHPdFWOZvt0A/SZqP7UqUWTIqgA5Ww+NfDyOG807Z7HKS0acB96RNO9csm8
wprreF/LrNYRNM6ZZIG5Kmq+T5PSmDYynBA7Hiew/Cltwvh/WiEtgFYy/WQq1qRlHPlX7PkqqeAQ
3pNnjYYdiiavut3qHUWiuie6wGY1Xbmopi1JuGPWOOFBiqgb7Y82uzuWbGPLAo7Tj8j//lO+yd3s
1F3fE2yrmH+6g5hQx84b3Vpyv4PR3r+uGDtEuhv4Zibvecv6SYqh4Re0anmvA4ni53sxMvkrfH0M
bBMBSeAf9ib2KkIdVVMx7AiTyLpvAnVgBnYa3xKo7YlYmn2Zuds/0WzMEdEZ/RKoYssO53yENjTg
mabejxwqXyajpNXShiGh5cMFNJuA5PHUGB6IBh1ka/Uqb4hplUc+XE0xiusLfb8l4be3JuHgou/6
F2uoPg2JvOB77/jgITLV7QyjKJkpUeOj5jq268yOcXU1bgqwcFt7BcOoHw4xpL/ZEUlVp3YkgcTo
zgzVX5oRLR/2jJ6n/ZGMzZLvUxKj1smiAcVKe+t0q5wDco+NM056DdKh/guH3bZFRvHXkdVdyKUK
7OZDzAK6zGleJk0x57WvYJHcasumMq2aYJs64OqQ1QG4FqWLnCgRhl36DHm3j/T9mkOfSJxZzgX5
Q9NlW2Ei9oSpDYcu4HwoI7+op7cADFIlz5rreCI0G2U0pEe2JZWDTHRqWmSLyH+2cyE1EFlLRRbk
GfXzwl5jJqehALchV2I5gDE4mYXUYC2neGQVT38iPPMpzwQ5E/Jd5hckOKtvvsfPEffQZfSr+UWO
hD2rxZAE9jBeE8SifjIlIrplsmpC92svk9v4hgKpnPgaF5/B6emeIQRcLMtrUVCOXyszam3jzOWE
kxihiAEl3IAKJnupnxRK+okblsCeg9rC5pA0llQBLyjQ3KFNCefHlXmflSyh9qF58CK1p5QSRnGg
UGlE3kRRQ5Y40IVHZL07pmTqj7BVVzyltoclHUDV5iMsz4v8aJbajZJiuvp3o7khCtP1mkUHAEoC
dhZIzB8u4sJ2Ysu6/q6kyxphaDkRIIPNlAbki2CDmpMIY/mZQqjbawWEulQupjbHylncLL17Bi3c
joVa/hvIGrEL3vU5UBwR3eIII0HM3UbWiBwBjFSj7tHXcpWITnL0LVRM6LYH2Hgw+h9OUI+HrJu0
x7BxiLUOD3zn/zdPju2EoPiBEt8WKarGJAhRDpiDClSyZS6JeDobXpvk3J0BONWSO/U190PXon5x
uguJb3PHwRWT8FeOr0bu1ta4Auk3VsJJvAK6xiKlyNhPUP/WI0iRyeyUnQ1XJrM1rLjQDYnRBgta
U38SF0R7+q5h8MG6FyDs1jPzOhNcZfTsSWPHs5dfHtwv0aC95kYFD8SDcu6EhqjnSvh+UtgyVec7
4ogxkGo9JmNRj/K8qLJtUklAUBzKMD0Wd18wDZircNFgDtpXTnsEy7SXiQnAP22dB8azb6Juuegr
PAK2t+BbCq74/aroF69f8cYS1IJORkm95u4I315cQckxR4gQkRdr2i5kLX/iEIVfrpMWWQGZfAOU
G6hfhgazxV3edFGxhbrUoUv2zv98mnvHcWx/ooDISIUVDjtJrtDUUF/qPFZDjULRzgg2RTG91kX4
B+MhvCwIFUBstQaBaRlA3ncAQ1l7ayeDgXmGHzN8ibuSfq2CQRMWBmzttxtArv00EpLBF6LxYEBP
n/qv/8vVrdT7ZC3/ChJHeO03WqvDUGrbZY/x3Zbm5sVE8jRuSshc8QeQnn6aoF0eQof9geqNOaG1
lzRZ7/j0MrIXs+KeAU9luvdnT+rRIE5aGuD1OGE2u/i0tVDk3d5Itf8Vfic/Dh4u254kHnlKyWJz
V0AhW4k6csw5sCYQUVTkOqNN22ou82K5P/6jrKEpOJ7+glXlAxCjhh0H8snNsZNAlj9ONiiJowuO
q1J9GN2/k1OxXOfMTSZaDx3+GMpwYcSqZTSAby0XjI/bYg1cr4nNTcMazJKQP+TQQ6dlSV2YyVIZ
Gzu6vWfeMA9SCECvL+ej/kzeJsdUJFiEU50JnSYqbcfXBPkTi1V0Xo/zTVuKozsiyhcxt7fIp/IF
P8K8W1YtZ9RpnDysW4ekaKEhkuO/aFl4t2TGhREejytkOxvspmLnkE8/lhl9jxJU9/X0nUDI5d/G
+L06xwZbwbJEEbT2TP9Ppgyr8hQDt0P5SGGVEFDJMw6123WuGU2a4fPsqaQrijiKRXDrz/Sq9mhN
1SgQsqHoKatfgJ/krtLccHH/4P2LbHKt+JbKXxOsFWRdIr1UCpe3nJDj7BMzRf9QWpoftrKgkKYZ
UrAqPyYqgwfczkhVLTTQ79hy2kqoHzPcygMdYO3NcPTVJzPANH0B8JWkhrUErtlmmAghYayRSf/f
TjQ37I4WyT87hF0N6FLyJSIZwvZnVymvN1QrNURelS9so1gH8PQYG/QNrZdx1Peno0q+oXmq3Slq
+qYblZ/ym7+Wvk8Jz2U3hZcUKLkvTBngpklOmrdbx+frrcWLYeMRTIAfnsuDRpG2OhDfi+0IFOUd
zFSO3BiwKvDeo0LN3Rt1B/ptpUwJ6d8Jbe4oU/2WM97qmG5W+7LKvLwc0vTBCIAh0YZQ87+RlPsI
Vc6LK4aWmZpqgLhuavlH2twD/aebl7J4iWABkYf0nYiTKTyHmBbX5zBrpbz4wk8ihAeK3v8enj2s
EhqgM7DwrHqUbh44db8TL0l3Fhc/f96kN900DE3otB7rzLmcrsW1TaqKu3j6+B4yG6wHu38BeiOn
wWg19XUNtnM3HSircXi2p2ec+GtHBU/yHpV4yUdXl4TwHjbvtzYFlhxDyib6HMMWYT+/yoNatXgU
F+AqEAOz3P7sqbmlkMRhE3aJsnxXghJPS+kWLqRktQgX6j1u6zMlFaliwDaQJGUvByW5udMvQcJQ
uSGMy5WJlfXrOI1Y4bUCrPqBtw+6lJg7ywxgQ0BlHCV0NNlyRQR871O9HpTmJ4iUbchOXG224ycn
g0Gvb9sNk8QhxuBICSysHEuZqJMCprYNFEO98CIXYPPRFcxFlwGuQ5R/jSXJ+d0tAs5sdA6VCq5d
pFYvgDRrgBBGiscCtYBs+a3sXDJcqrA8b14ODO2vUwh3F4jOBQ22AOqs8GMORYOnLic+zSZ7baMT
5wTIwv44FBEeUkw5/JEBYN0nye+oVutOCeN+fYxhjWiPlXEbQTWLT3Rlro4uDf2NjxtuSefGMCVR
fnvhqSy2zBF3tV9hdbpaDPNzoPfZ40RyBfRhbw+B093GvL7pcd2jNGQKkcr8VGCtI/Zun1nZ2AbR
9UA35Oqj4ivsvL75sqIiPOhKpq+J0pKfIkp7ptGeFpaayBVeKMwUv6QO2Fu2LbYqgWJsdOZ0zbwd
+Z9FVij7iIATgZEiQMGYA4yEYcNCsVXjWSUn8d86UQaB5Q95BienzhF3p9LjvMkSfGu/eHV/ySIf
bCfCeJuc8PC1nVle4T/he0+REdnSLxZBD5+h+Vf70cYgpwtqscncx/m3r8PASOH+WuSpR66gnRL+
6XygC/CuJWnfwXqTPGmrD3ZqD/US002A0CsMS76XWzpDuOfdyze2E2ly4hHo1MfE2yE/lpEDIkko
U0LW34tPqUJvr6zDAECSn4PlrMhsOdsOvZ25MZvaptCGNAsz63s+N3FwxpaiB6UaeavQr2QpYevY
6H+cM6c3456ZvLGrNh9i0h7jQOnDZHoHGfnTMkAyz+iNm1/2sIrwdqnRhELg5l1dJvLEcmg1LCZL
neoF+ViczBumWLU8ctiYQjvLl4exqrwONjbYL7xVCbHJxHwBWGZHz8xlDOEM4zRluO+pMjb+4DTV
dFv/2Cc0TenLEu7ldm4xZaqqCPDw1AtI3s6503uPSZtD8G24E4kpu08FBst5WnM8Z9Eel3Gs9v+u
7an77RcG1MPoZbF7qu79htqoDu9dUQ8qqUmIpE66sveah4utsJatsIJyzL/HFESNuW6U1p3ynYdO
XMulAf3+m94q/jd8o9gqknMo+Cd70Y+iMPkcUsVozn5JCK6ldd+RXGh+MUSPQx3T01/uwStOEHKB
UBurOsqSmluvL9i85piQBBDsuKiu3pSLa/tIkvM03+JTGlr7KHO1n3LtBc/2cdwPidSsxxL9PTwX
QYsc/Vu6W+AlfOV4tNfqESkmx1UIIzenFD0eCDyQCuU/uMFJyYmrinMJhXO+FXZYNYVhtN2/vAju
pslnUQR7KwgJ3MTWRYtJWLYZ8hN84JDFth1hXRn+2cBk/f3kKoWWv2vYC5VhUsYl9uqzgZ+pKK9/
rS7G1JV6UZGNvaXppCvssWN68FG02y6JyItTi8hX4CehuZm3WLn+PPuVzssRinMD7kSoS3+4+sD4
2mQ3d0LN3pva9ggewnX4DMyx0UsJUF/o0DG6ooiYw1V7fHYkrBApnhRax7Ki5KPIFksJYN2qmYv9
MiA0hVG/iOk41qgJF7VCchrz4lbJc1SaMU6g5xdM5Odit5/N3+/PGBHUZCQWZDAKGdGpT7wmLlDw
C15q2bKhHLBft/GXM8JousJsP/eJZe+Cx4tZLqY5pjZ8qN1ojbsbLKGYusXxV/TJOeiW2rdmPlwy
49r0C90U2rT726yLtOxbGcwNLzURypGBSpggYUORhPZFdSfAI+1fZgFrW+LWw8Jl9c2mfH5PoIB2
3kOG3fr0/6gQPis+eHpagl6die6U8Dr2emtHzIJ8IwVSzkxhclNKHS4abmjNJoDjPoAwrOMo1e+I
lLcKUlN5QR6iG9FbhhjBKdWUsQ1L5V3vBTQQTDL8POIfUOWb+Sr1YJ/l9FjgQ3jRNZ29VreJvKs0
i6tB7KmULy4SqPCMoyjiv3dDoMJCxL9g7O+br9Z9KICywPBaBLxJNd0nFExhORjFCGFd+DN1cZmx
DAjokZGnqL6MBrXWiHpZi06qbCFpgOfHASBVEkhtuSdfzK+caSqY1oYzLehX4DE9sPOpNhvO8bkp
gRqQlOVxb8YyQD5+0RjzfIMpSERDKlDaaiJ/+LAt76D8MFVaE1i/+s7a14xaV6KpeexrZnfgfSZi
8IUy0AiQFlr5EGV9YHhJTw9RLmTJHfH76RWOZ0YxKPTGltNERN7cg9debc2W6rcdmWiiEyrFE0Zt
CrRQKouFBlyPPLEO506mCt/sKLZn37Wqj9eKIV6aA1/2HJQlul+evTRf/AMc9ueGET9t2YbyX3kJ
uIZjHTTZMJPesnP8DaUEAxrqx4kMW9jUjzXHKKgMS6iH+bwONpWlot+cg22fW1pPHw7vs0R1ilcs
wc/SzjihodBhpTa24xDRnIuCVcdM2QrczzVA+8p+Fk8Xk1mwt50IH265hm8lAGVXyk0vk8SIWkrN
+yy0+EnvBdun26tl7phtW56d/LXOn736cAAEOv06vuh3GMsOUdue3bChTKUI9+zvaiSAYJO4X0nt
FsRVycHgu8QBLcGXMsLgE4cIgroidMbjEevG7/RoQqU4CbnvgN0CgR/IpI/nvVcXjJ1T9leaMJwI
I32KNWpy3u69fAbTjgwl4A9WPQkofUguICqXcMqgISrkqJcbiErIcFZ3oMoOwV4nPsgxZj5wY5Ho
G2X8vke4a0zYjP0fkYEzrLdG8IRbD9fRQZB5iYRmOxed18O77W615cHZmflUD5ikACL1EkIakph5
JXqRcbyTOR6u7Se72EWwrM2JBhoeKIpGdbjsnR5sQaVMIZpywkJxoIY2V8/jj11egQb7jmjuo/SW
5YPOEIfv/MC+DUffdCPRZU7M68v15vxfqwdkRyLJ+fUkyBRmIN/R2/2NVmrVunZ9MU1CYVeV+77e
gR/PTuxFLCCdc1+i0tcmmrkqixAw0dUKG+T08r+YLwz4lgBE9CulL2UGZorTNkNPyuMstz9JMD7c
3uPoCsOBh/Sd2ANqAQw0ekSbPU61v6hJII/VW3S20Aqlg3XmktctepRLWY11jcHYM0r+59vOV2Ms
Vg4Vs5pyBIZU8J5+o1enwErrrF42NVLoXw093HUKEwAYtWvP0qkEQ9XR+rYoX14icXEn7fp12h4c
vogPjlfqZc+DOIQJqFIkSqyE3Xfd0/5QU/yqZQXau1kBLD7xsAZxOauy6lBT6OQSUHAk9fHoVaXt
mo5jh7bZ6Jl0HeiSYDcqrAZDIzmoLt2T9diC9DNSgL2JtutBUQvNpZRtZuRSjLVYhW2Vt4afC7Hz
uakNlmMv4uAi1ZFz7z6W9eASJx3UOVUAPTzZSzyXkhCCq6MYPUZVXZMd+yC4AuxTkaiff2k7WNAq
u4631vtCiChJZCpHDHqlDZ/WO5bf9kNg739EFaCtZqRoZtOJXM+BzIH6Az1jP5zWDmrmIzVxJf1l
yu/V/jCxxh2LlQtz6Bj6nQhPQzE1C43sGtXf30o619nhkWK6Jw92EgSGxMfpJk4KnjmBEHnCpFYI
8P6JIbj6aAvB+jbs5nnLZmbqjelqkBhK8Hdqhss61fDmjP6c06XTQx/X2uzjLipmlaTCuUVQwv+f
vdCLhAP6PMXDeuag4Wwzfo/xsxP1c5aSzHoHC9J4h4j1vTlBJ7RbMQUEa7nP5PHtULGkO9lRF02n
S6OlLgvRDEprVrMoCSIxIlG0LTcklihbN91z1bXZEix7RXd5z6iT2EISZomv9e35+ADVUpZM8KXK
Ye1LYux1fVfpdD8yU2vwTnmY3tWOWHSdPSp9af2vDeJGpShAsYJbdDSCQdI/PGXBOOTLNUnbcnfg
o+i73b/xC2A6nu0VZgmmo3SEb0y1NU5Y5gMTqlYwbYb3L4gHN2Lgjc9DbAtM7CW56geGUBO8TBqU
1MnHJtycKrQ7ggG89AS02zNeqZz4As7XFOBZt8shxszqGTemXG8jwWeG5hNuiFVtkgmPbE+iXza/
M2TT9rVEfBZYCMUgEAGnoy7YIkQwMPSYnOl5fAiuEld1dRdPDaoWqUOD6JOVFIye4ra+cfEksrhJ
EHNHYoMcJfNxfggB6EkG1uhfjm1lFhg4xNEn7e0u6xQQc2t3tpix4TMZX7FiXzaiOxvd20Bu5qeP
8bjn4bknN+48Dn7cV1nYKAj1GNhAeSeCDNhRHWeqSszy07kICzbbwlBGmOn10+yuvY6TG86Caozo
Oo+C3gFNuINdGsgQ5Z6TeyhayyYRVLZUIrub/t9oJ32ayOjlNXMprkFGE29ERmya2BMuaP69rum+
fyJDW0UF64iaI2gE1tRYv6C2EHpXVNOHWvAjzy2xwOox8SrIsx5WYZoh+APp5PfFfaOC1C+WAKrh
8rwnnhlXnlmP6qm55IsaEZ+mKU1qgaZcIZDUd7nsIVSd4XuFxjjpJiLQCYuSBCayKiZWxKEhgxGa
quwFfSi1AYc8dqn2ZcZSjUopG0HZiidLb2ERVJ/QCdrLDfdiOBi0nuZ1iz8gYWdClDZDAM+XlFJP
AhggV6g2P2DjpbNPBVNmR4WXslikDvKuM3vsbkcpeMhZASXNvOkA+Fz5TBJOqKoHi9IGCnI1h7yY
vhOjMsa+qkUX5gOHFwacdUfZkP7ZAUi4llGEEYX07CgwZ65edXcZDavQas3wsbDgpbWkx63KVEtF
p03p1mvHtdOuaxO2Yk721xWtN5xY67mjo8m5gDFLfVn1DmnRlF3JG3CUGGGu/WAXDhfkPsYMKV1y
wC4UdSyli7R8GpUe5wInc69gFYGkCWXRcmC3TI4HRMWRKw8srvHlzYtU85+BsmPx1ZHVzJbm97Jl
I7unEP//wIrqrO0rcRIZYiWZ5L5KLftLAm/OLzAbCnds0D11Ugejd4SOkEl1Q8bqPZvvSmQWddRp
4ZQ0rsr129lhoyRNAPILkA02QJXUO2d0VK4IxtsQef0Em8C17OMl0APWBMR7baRJtZyMBjg2P3IC
SKVcr5OiL3yHMuN0U3SHxOvkVJjtQwfQd79gqXJPZdzLaHAXEXyU4qmTxGfIatS++UD1ZZxk6hdi
14pYahr8wmjhA+1P+04eIxFAHUxAXcQsqBYvlMV5bIg2hudKdrsI+z5j+IAUM/xv9cIHvcBq19PX
IJUSh1EGGMpgQ2vRPuep7EChxc6AKGRH2agppB0UFQPrCzj8D5ildsKEctDhnsbiv0lC2GFYxokq
f5jBgC7pYIJKAZ2JZMNQMenpglE/zLPbh6qNdDxYcux0MfcKCEkXmm+DnkO7ez18NtivomK8VSNE
6d7hAAdPcAVRWLIF5iWrOZ37Rz4U2yRlCv+YKhTBcgMGlt9DRgnpNk1pBfsLL8ktzxQMJ0/5enFl
eMNUtZHjD2FoUEzlWiIJHEceoQvEnQ8OFl9jc4E2JfgbRQguUKMJS5mTEsGSs5V26T6o1aFaoNK0
nHKRA7okZcsCZxjwpUf0/PXxKak3YMNQbEEMe9tMi4zt7f6+vp57pV6U0eZTPIHT5DLxfLpXkp2u
rqzI0jypfa/VlzU4Rl5jcpnfPXsxjxM+kWKykDb7wQOOy621wbeXDnwHUQAJIkTl5ngDW3sGEFU+
Bgrs8P3AAMd1kNY6TEmiNeNVVR87NRmzA+BhA7WslxyuCTJKcEUlQMtwMtSRqQq/pubTZhmDq9NN
el1S1SF9X4TO03EQC5kTvMPs7DYJLaRcyEoqdw9amJEsKKpH1TehpmOwUHZ0fUh8UqaPe7k/UN/L
QXrwYiTjKUadSIkWFP7LmqqWfUy806qICHuZWMaEbl0Q2GwmK/YijJx8KvXb7Ypcu15d/C/o+LFB
py+v7XiuJVYXmvcTVxEd5Gxm/ZZJNJnu3rbbKE83q61e5ggJgbzar5wkRcOiM6+Gx81WKYQDElAq
6xswO318qfMmduWD01HvFA3DwnrpcdYAvfVsC4xajzJaIX2bf3es/XxpNpYJci8jIRdwsQ060FXk
rPC+yebakj7MfNaI1qMwPh/sRZgVY9gDLXnQSaQjGOx9ZVRaeq30gfB3xvxpS6jXxRxHclvOH6eZ
Erm9u6a2Y+L1JqHpXa9LZZE34s/Ei7pc9dYz+Fz+2dAdVQ0iurm0PmM7OAyIudHnYeYAXrG7Aq2d
Eu2gEiWDaSLRoQOWv8rF3XekgBNxTsry/NO758J29Ump/vamXaUea5svfViXDVfqLoEivR1kX33W
LsXk5ssyPvWxnBBKYTFIcDpxqJSUvRdPGbbXP7xBM9OeP4Ew3jVEYQ+8Mbo0ZpUmtR3q9dwJJ+RB
VcEe2vMEMsdxlS9Fs3PhMsvu3KXMyn437Dy6OzJy9EbFaYEU8q7d8hNJVaDIVB/loOVkut2S8TkQ
/Flw/ZadYXomFdpBjS1uL/L3LFXDi/oZUlaKLVMgN6HHtj8iR4o/tJB/RG8EP5+PKqP0giXv3X1s
+gTitjTbnWuBTksPpp6V6ywG0Pw0HpPShymgv2Htofcd9Ym5Zvo+VYUQlfqL9s+qi5UDZYnvFWVE
kHDdRyRKkMlGP9m8GBSjWpz+Fw12+IL3aGjyCiVSK64eHhNkmm5d41dCDsymrtx7GOSblg3NMfHR
PE0mDbq/uaInBNa+3jL/FotjqV3hnDaTPIXQJ71pFqnc3dIJSHjkyQCyVuBq5l8+Z1tvo/fAyxUX
UufbNUO0yBlPCyTOCSMZYblewH8b18jAA2NendKvxyY8LQpzGcjEeuHUdSeke8HEsiRMUuN1WpIC
3mKg8VMlpPjEFFgGJQOjk+NcCfQpu4+0YKouKS3xd5BXNHFisDwGbT2cspE0o49iywIOpOMlHj8J
tfXEGFBRmqW5nlSkpSAxCIEOixJwKfZg+7M1uD2E4hfjGrYkpjjyFwxeR7QfUhP6yyQgmSsSayqe
B8HBIGkaibpm8urOm9mfnIl7/eY77m2JmOwCQRo+LoCVsQ3XlNB2raqRjlnnwXM09B+mh9EWHxSh
fxAPikxpEvuq/iPaxPZ9vdKJqSFvovLyubaJvW8Ki8j+JO2iy8COSt91U/F6Jvo9Im0mqNSibTBo
0OgKGXQ/Nyx8aCHapRlY8FhdBq4SfsTej52d/lPJhcQpwx47s3+wSAl/U9zn06E+761fHdrYtgXH
nQvoU1CfbPkvBE7cX6ixJYeHy6n31GJkaILfsAacBlFjXl2xjkR203t68pErAEIFKmFKKdquedvK
lRixrsqH9bXHdPGlTkT6kTQripTvWOw6ux+9PpjsvEaqFPvPnsC0dRN2bUiBxaDNhNekJfM+cHmV
Ggod0dSPoLoni3MYh+IunR7n1RS+w5ExUmKixZNWnhGYkbq6SWGDAuGp2BF1AU7O87XiBJp+vwbB
k+Pv9fhCCJ46vrWuymYqHAioKpXo4tWrPXvWjLOMFRdj3TDU7KsCoQsPIu6QJ3DEYg0qSP6MZo0g
7JR5NJ14g2mB5HOvr8Vcos9CROocxtj8kA37o5zchaZgJDsY+Y3rOinek46F24gdO494K8QRRbNe
aCZ6F39SZ1p4Hbk2q/pTX9frq2ydXhFsqSHZTGeAj8KWMYcb4vDOg7S5DRzLO7hf325y5Iuh3ZRg
xX/bPHJkjh5l7azumUDZEMvfcOfd0DVbM47MrDaU1KXV3+6dpUF/4zbrLZ23inFX4/TNGmdwViH4
LnQvkiU3g71JJvz9XVFxuW/j9VcVf7OfuvaGwveCCOomFeO28WZBBsraz6kzz2nDzCleZqoAk9IN
bAEbfHB4ogogh6ZTc3wmFUSKdENsRmfCL5DCeO5HKBQ3zYwhb//ArEl7ekOF4eLAe+Fe00s3qqC8
U0WNQ9rVyneRhjKrK9/jmU5hOL+ovaGYmbNTcEHOjxxNOQ0italEshKhwvedFunEV7sLY4xe/COj
JUpicIUI3F14d+qnlvx7LWwP0YrV7YRjJkVRnM34d4Kgs7xe9AZGV7JuGzxl1BpufjlLECcFAnOu
202BOnbFzQ+nZFMIrkF8/jYmPF2ThQ5gcLeo7vDXAMfvLP1wUgJ/YSDxo/3PfjD/7J7iu8dtLtQE
SK//BETTgQ/LIOepQhRcTTeBdsSwgucZNTHgOeO46Qzy6wmVgt19a2yeVEY7/SD2UAUm9zZh9OqA
tKJBIN2DJ9ipzbZLk4urayYj9TLIaM4aPQ3qRdco7LP66APy6A6GrOVfEDNn3jtq0OauhPJqUIHw
xO5AO5xMaKnrnt4jM0m+GZJrRJqmBBx8KghteZNqXDrMF74++wUQu3Xu5zQC2XR+tVeIDADbGMO0
BcCO33QRQMJm4lrYgUqFwkdmPUmc3qWQRXiMCGxeWt13MTooH8/i52DXdY02msHnEnJL9rb/94zY
v+D7ocEJ9DMzduRQdUqgpeQgg9NzgOz3oHu4ZUah7VXqusk30bhMPgez2UjTWEKGBVwepRHPcylx
//qdd9R8D8dKBqU8f5MxrkrTFEw/bpdPWI+VT0ZfcrhTn1nuXzlcfqabmHv7hCNu1HLfuDhQuPey
2dkO+UCpsOZW6R8NOwGsIvHI7UJsjXKL51uZbh9Ti4mXQPkIpgfJLocFFrCCxoSRlKlrN6vJwQ/j
Vct0uEDTBvvt0FN6UZYTnRSr3qYKBuTPmRDt6H5W2VQ3XYxi6/aEFa08LJ15h3xTQ5LAVjlfSwzU
GR+vGO2xq++bkinqE3yjSW1h7pxV1VjuACgyt8qSQJ2bgUh0d3D7ihByUPVlDdeHRJVi44aYOP3P
lsCGgb8eeTl9SmeEFVQgrcsXksJbrXEtWnLCq++7fhUT8/7sdj9CoFrSlKwKm11NjT9rOTJQuoOg
KvloRXJN485h1ZQbnrtwyUgsah1eNMkeXzOSZHuP5K7EEdHxYqZTGeisEDowdPpcLqitdwJjYHlm
sUR7kgYVp6brUeumF+S6ReejL+SIjDj9AgIfa8Wme2ulMq91YYKje4Vp630xIGgNouiE7OpEKcjL
tJspiEIWqtth13eSiLvvjJkZZIIfMXXW+982Vtp4mAIwc2bWIavgeGaY0Iih6wY1tBD5qNHJAHT0
mRMpPG0vS3QdDz8GLfeplUF1DWiwlRWyltZRO79IX5dcmAcpT6H0Uw8OZVZir4CSqrdel1fF2POM
HCLDTXJ5EaksfriCEZ/KHD0EH04imOYxeZ3Pk81PoBrcKKAEzGOOsNyErpnUoiV7L9Bw8DPU+1U4
PD1btivqfU2c4vKVnHWl1JR0oWMrnGmQWRLHSITk/OKzcE1WErM83a+H4vVDlOGdEP1SJq4EQV4r
bCXUZKbxuK3LjjpLotMRtzw/1ttkQkAdoWsLFR+7pcucVFPi10jKKy0GZ7WruOz8NuH4NycRw19t
iOL3TPjZJ3PZsJJWT5TUPNtlY5mw2otpbFxIAh4GX9+m2zZh2FFtHv4go6YKm7XJuLt0bOMqFaR2
Xr8JQoQ2xTm9V5PW9A3ndfnJ58y9RA5ELeSGm01vzmtLLWBd/KIM5t37mGseskO5BcrFM1mzTU3x
H9/DZ6TU3ffHocbkRZvIlA6IUb2UQwSjSd7CnJwfjr/Lm4tBMjZmfZ7OQdVqfPelaWhoNrP7FpIK
Ezm1KA9ik18BVpdemTK+ULRNKpQkNx4vOTR39/mm5e5e30eCJUU2zEsB8vAtjwMwgM4xJWS0lZvM
2W6BamiflwYTytqiQZAxC4IOWTHUwM9cHeMIk5fohUY5A+sMqcX33mV7ogdl0+vDOi0RwJ51wjO/
z1IjXn3MTip+QNwyakZmt9ansWLOpGlzczlRDSDsB/jZZmr9JGD/8afcZwKjmGTxIltoZT7EgcNa
uxXVg9tXW7+cipvwxXt9vCrkTHpc0mxen+rxvArBWyT60IW0tj0xyOmfbufLYxmPHe0ElDWC7uo9
Yx5uBemyCbGfmfcI2YNIvQTQxKK7ZLpORsbLPds2r1Lfe+Mbk+f9SjatbSTk5mm5QmXj2izogDMi
7kChZqQzT+vLoele1EsZM3qn8hcnclkroRMNCgTXweACqzXV482T2YdxqIz/hLuCCPMnhTQx+4Qf
+zGmbJ0VqTsf94fFXJxYozweTk8k3/Y81QPBP8xl8cNpGeZNpx1ecw3hBgdoI1GlRRIMyfahyOn2
5Mz0n9rl5Y3ccW9KGcwk9aZsB8WvSJ8tVXmUctEBJORMJSb3sIYKJsBljmQJSLUROvi8i2135nQE
8wiEpgCk6lm0dY3B00LTYsXUYfc/cyW9lRg2vWUReEeQMzUWgt13qSSwQt/ZjXpXAEqTP0H2MBKm
+3MNZbpjmsnxKRVtDmQ9lZQ0XMqn4ByDY+WnAtjueJA9zE/LVcY46H0Vpe3+utW3c4chd7XC567H
EjYBszhQ+x4AKQLkj11jemImZd8Nw0SDGobcTapV6uDDMv+Q6EyemVTAAlUclNRAYp0/8WwLJAIl
/Qw8ltNhyzVb6D2lYSpN00jI1c8uzQhZKlHlsDz8xyazmVLiMODPRyS4GEzSvZSFUPmkPAuGyyVi
5Vcz+Gc3Ux5P87dwVSUED4nmE9Bv3ys+93enPefNyfV8h8WKwqLapXq1pK3RibzE4lcENmT3mKai
/79ofIMMq1jRhUfCIUrOH7qREEtMIe2KGVPJSSDdZ6xJo6V48eRpVWIRPL6U5n0+iTw2d0xtxZ/J
B9H64kqr9JQAaQiyjf+nDkuvnYpnaX7PebALzxwH5vKeqGyaMLXXTdcR0TeIWmhBRZaCLTioNBOD
VSURon7axFoPqTFlS0MybDNkSNBzzIgSkEgZyiaUrsPxm+gp77uQ6/fL8S6s1zp9+hU48O/+nVHm
W7w8DN5alymWwxkxUU17XLghPce/XMFT1UfcCrk0cVuktt6SKE4NF1QRlp+zqfEIPEGDDiP2E0xE
HlTt1htliNvRFskIkFs1yK5xaGWxgZVujF/XIwRNOFa77rwKlaBRYwrPAj8fbe8STMlQpIwuH72g
unHz5MPA7xJTgMHZGieTQyoTR90rIR+wWjzGxG+KbvZoLSIPwAkevUsG/2zbp0h+rDoiidSL0Mb8
xojZkowtXklvV3y3kPvnA3plFBFAFD0vaG3lxg/QrTW2p7DN8sytgOo1bCVwhsKSscn4IQplCrj5
u53e6/pT1z+0vAy1aSQPj6iL3Wj10iYS8EwLYUi1Bh5J1DwdZ0VR4w2GGPheS/99UJfRXqOUepD+
/+tdD2j7r58nQZ6fyAu9X0ZqKmn+fUf1RbG+4P55l8WcNyAQbFw+JS9wpeIMpCygDjlyXKpBKqHN
PETu5LM2+ku6rX1+jqrIweDG5HpmPAbPar5XmTNvgMBKhK16qyhfdlLIkBl6FzpAX5P3TyvqG+rO
YbhjfIQod93HT9EIcmyqawAUzLSfzPo8S9fiSuYTxObFFSXhwmGXHfW5fF3Dk9MUNLTj+NGRjRpy
D52DlVbhdUJsT7ffpVeuKGQ9WA9byEWs3tVNRsNHHvTW7GloCEZe0cOMcXuL1zwuy048CZtjvwoS
X5Fot32UpdBeH/knscSC2TC+XJnJas94ZzhfXJr+lBUjaSHBvpELlmMQT/zg/DjPWdzHUp89vHbc
s+Q30OFo/456mw5SCXx12qAU36mYFljiS4nR4Hye4ltCVTzMRQn8MRXqHLkf1pCCQpFs5bc3ImNG
RQ8L1YOfhmoemxJAFf/3C4xKryubhZv49dXyfJoxTN222a9zqGo9TQsjFUcaED6I4pyknV0ujzVj
kWUsQnM02ECDyF58hz2ePPHRPgoPRY3Sc+0Mu2eNgrguKI0fEArPhZeRZEzK/wdmXhU6UE3ld6vD
/xA3b1uxN43u+c1wZyM+Y5NTnyiJ7R9fo4/L0g3XY817yIPntRBl7CuYND847FSXbiq+Mwn8D0rE
N+NkMRwk9GSQTAg6HvF0kneWLsBcKouzyn6X63MHig+UD1ftzt+QLN0edMMflg/nRh3FGRTfWS4d
Hmpg+mtLjF2MvniUIXRzTpINwKVq1RO0dgbWc7PHj33w85tDLU6Sqvy5W+Yh3TEHEYef6Zyu2yR7
jjdV2cRTqJarsJ7AbiuX2jwUYFuVwqBzQ4HUIUugbnpV2nQ1M3WdT2bu45ApclU69Td4tPMNbLo+
yYKy1CWtOmVnEMGyLVwPMlIaVAPhWnxjYh+Boz8GWBp5tghMSl6gjPwL7dB33H69yzF0gplaeDS5
SPsdivai1ctdeWcAfeLp07KUVL8wS7HuPbWvZSQ8ByTLaorfWbV71oHC30VustQde0hNr6Xq9AOM
5XmPMfXENUIGx06JhshpcGpFkzhcyBITOnL0tzFYN6NVGjRaX2rvaBBfKCEYvHmRWsG2MiutQ38p
Tih+oFMQbpoZ+xuXImIYm507KuCyOUG4nMVCe2gswo+KWRoDRlq2dx6BbBAxVA8x4gUI0q2khyvr
6LPq9lEHu7KlyGv7VYdBUAZW2MrObTNM/XZ7zRT9KhmVSgoRcCSb188ifRuwOLQmRcWz9bt0nJXt
xqJ30gJu2whgjbC5/jH+d5FWAX97XPbMVBp18e0MlsLRNuHuXLlnHt8283jJOTEqBaoR/oA6IMBC
YunQg3XqjvnQbJSmCN6RyJB1SjHIBFN+Y7Y20FTS8dadSx6sxyCsYqNKf52NalowU2vH9/ejn8sw
9SkbLG37E9bCcfY/TBhq/kFgf1ZNMGmU0Lh0DZOnYy5zvtJN2NThPAHa2YeBRHsYUI33m7SyMCBy
p9eKHY3hUe3LvPdVt8LCm7yFqsU8vhIaxjrfJK2uYw9dzrjEcJ1/ucVNjAVEUhytWAcKk6n1IBmb
EzwJ4OMSGoexU5ZPaDPWJoKDmllwXW3nCaalb1aW/FHe+r2H4RxlXNJv+FDQX6GXXfp2uBuvDoZa
Tc/tOaWx1vV0DnEnNOrqazFn4fpbhmTssx86NZUGWSHr9ZAPVt66L8AvZMGy5/5hjG+V0/PX29Md
h0eS8qZur9dZcVA7mC9EF9+TeRoJXcKnolR6+tzsT4M9soSDwwg4BhCl1dvbay/mzGTsHVIFEn4m
ffQoBta3BdwuKSH+VjkrURvphrlyHNIz8sENngwVLwY2U69EhCSA79RKfwb0gbg5I01QPhu0wjbi
1BPI30m0qvPc9OhK8/+rzgXkkOJMSgWHc9r6WilDS9JFGaN2VOg9tNiQdPUfnyS0TamChjCL4dTG
l1M1ezFyDjYLjmc6A63Vl9x3l8lMalmF8k/bLdDWKC7tWfI1+NvWKMuO/07378Ef/ERvy6fk8fp9
DnxHqEMw+fLS36TsP62p+HtLItxuuQxLif4tOzehH5AtCzIjgidRKYP1Niv1TVn0ursxLqBiYtc9
J3YlKDMPMMg9fE8gUVfRCYE//GTm03OZLoUOmHTwNlXSnvToHkNS64P/MrPD/+CrLiHc422NKn1N
1QWukVFl6ABeLeKEPka2rQi2vFDPs4Ot8oDrYZVSnX5iGe88XU3Yca0odWDQ3Zm9vWEwJEbCQfbm
lj3EEbyFxUgAVqH/6Fq6+HQQzoQZLejY2V7citP2kA/FBOgV/girpa7zhPJgN5xSTc8xblAJvLNS
2YpvaiNAt7RQodkM13gZRKapUBgX+yUNyFvlC1/Fwl8zb73BiiC18OqVejcu7kM0FWM686A0FAhM
ARgp9ffJOKgo1+NAWI38NlLd/GutncfdgZZtwgeVnHF1r9jVZQ+CqlGiDI9fX8d/ud278Wp0Fha7
U7+SaBNL9tOqEXaa6I5yne9tzjncOM1Z/ht9uNaiz41m8A8E6agGMeFvAkXrDNkr5FHFz8qQzZ5z
+EjvNVm/98ak7xbU/mSTjAJjG6UN+bTKq3nYc1Ao3GHvoiHrxTYyLRG165WG/pskttJkm4NN536I
kT+612yATzhSywdKza5KgCqxXdzPhxQpYdARC4QzcPOu0q7xOZl1iraEUzNfk3ziy4TPbJGcv7Fk
0AaGNpltR9KxW4CyQoPNhxBdTVjJscgfgTCjpirB90/KaaF8HD1nROgVhDK1A1LDbmVT28ehk08G
FwmMvT/HOYAf6Ctjz34XVvM6E9KwnX+Ug9TxsgBdwrE3yHoA6kaWjgG1tLbZ0E1UZC/ROccV01ok
wTsqP7jIOsEvTTFV7EHKkUMV/2X2K5ivS8hDPv5aVbay6ATWShaluEu2iZ8FmmI9l3QExl5bhrcu
Ze+56VuZcXVAgtIMn7KcB1fbrUH5/MV4IoGrmOI+sBshgJxbKoIjKMibi362Sq80E3eFc/4N8EyK
xhjcqoaDopKZGwEcUgzjxJMZoo68jJUq0Rww2JDkKfiEpfgNH+IwuG6ZD9wbbjUtmyXfSw/lj/X2
r9v2l8x1MN428JgylCrZ66Y4iGLKngQrHAybTqVYwdvdJrGWjdkqR2OfCQejvZSx4tx5to2vNa4V
BNK3QOh+DSCiXaCtGAFBA/fVsvwkyv2nZTkt91ekfst50R04geZZAj8XtqhPtoIGDxG4UVX4r1RX
iEHFdWdL16LcM7TwO+c8RnrWSNRIoz9BxeLSGM2NByRQzyCk2UiiLlPlJwFVZIR48F5btTj4ZhmD
Cj5mz66UpHjrqw4nCdxdrRAphrclD6QRXHTOC9ztRk2S3cAyn7pkvOXxNBMUtmzlzmX6tckRlu2I
/DAZq9hu4h8nqCobg5lJarJdplk4WBSdt4nmPKrm11zpPmeCM4HynoIgIwan8s4d5B/2zbeNee9C
z3ZAuvD9hQJ15cPGErLDQx7OYio0sfydIYMAki6LIhv42YopIk8o5qFHPOlO1qUoGqXiUmAH3vEi
41TKWYwlciz5vxBFg2cGLgZAJv0weK78aewXoIW4KiyJU1SSwnsq6ECRtdnSFl/Aqd/wnQKoQ4JR
0G9JMgUM5rU2S13baOTeLzhWDnSsFWOS5LFvT/LY2zKJWZTMHiyGX1tmh1Uj97zVyzijCZFd3nsV
ALavQ4RjvGQZ7bHPeDe2PYPP+wYEYCA5DmgV1/ERJSGeaq8My/QGjKuibMymFjOxdzuPAsPPetiV
2zuQl9hzLn2RqkJIi/O4DNKyeT0TUzygCxHLDZhVKQnhneP697cbfGzWuM9h2x2cYB0mOYIyCQGC
i2ENUhbAvTwo5FSQZpMVTaVgqxJg0fxAcWNcV9ttSG1J6fCVr11ce2F35HPhwu/lemhq35bFKbOX
y0iYqCFH4GgM0d27R3Rgq9hdTNzPE0SCJUCSJCk7U5CvoCW4mecbUHhAdI6AmVSFlZSMcXuqUF7H
5507/sdUXUNoQn0WjHu0+PA6zINVP8QtzB95BRs/PDfW60laNqii/WUnNl9mXzkotxa98iZRRY8b
5jY0XS8CTleHt0JI+2ZfW7ImfFFgajeEMWjRlyQbfVMquyfz7EmdM7mg9iRCUKk4sFyH8q3+b0np
OrhzGVzJDaEYPWz8v4p53rhLNY3GFRadP4bSvotzub3Fysd4ty8sCScvEaiWwUVR+0ooRatn0v4D
JIvYlKQL7TGr34pWkgUei8sR6amu9IIBIDAk+U1yAtxgofOOaboYa9FB7+lWFmBJte0JGBtG/lq1
Mk2+m0jzgBTNTr3HC3ogxR7pmzNmGLMTQYGqeIuZpCM6gpDzIWYgXB49qo2gfO0RiElHUtEOTVdp
eYHdYQ8jfLo87eWDXWsth+tAsXM1o46JcfwZV1haKVpsFbSd1kMtFmP7e0NuTwHtSq4HxSh7Ku6P
bSWwx+vo8cL9Gr1oQnkB0loR+8RKRRc0vqJ85muu0fkmlT0X6JZ0hKfi2QpznrH+XO4m//BGsgia
S7CwArhtP3W+KJKTQtWhcHWugJQn/GCvs/pdbg7KYbKCYiAQAc2kurHiXf6eupNj76MvK7T3pHYO
1FFU6Lw62H2NbmBiuhFlw02lUi1ZlqrKR9Hq2JXao/bVi22dUxyURQgeH2cpHVC6cJUiofhfoA5c
ue3Pt8cCdG4bTs9Ivo0qeJ7SRQWKwxrhp+1Ori5ZcrNPo4PBqMYNcZMjHvfSvHnc6epVUk+oXHyA
P5BRFM0V1ITUlNySqFPZINmXTIYicR1sevheTTpizQaBcafa0mtIsrUUx9qyDJrDwkTnpqAmoU22
NGzQ8FFvRfREl6lVYbUaoDKN4xm5a9U6Blv/e98T/ttFUoGnZx69mjllH3OZxhG1imY90Np7iRxn
aM8vQ+xhq7u55HsIeXf4iVPOPEYtd9QTFznEDWOVILvA4LEbffc4i5qLyw/w3E3ziGatd2x5XOqX
HlvH2msJoAuSfQOv3+wKZl6xk/2nJf++erY2EW5lhBytoPtQHgACc8Gole9kZct4hgnMAFLXfcin
wpJxsTXzY8Vg9/EToMRWj1z8QFJbSpxIsnZp/BobVHyBL79X06vOpj4BDBRAUN0HXL8ypZkCDhR0
2SgmlSNk12TqgUiV86dsJKcaNMFoebnPXn0ZOLvQ1i0133Fpgzcz1aKn6zvvBjtoLHYcDJk+M79c
GXl2kxP6noG4SGWD+FKEA8dOkG0BkMV5T9fHQDrpu5qzc9H3pc+0HFwqm73QxoAZ14U0s/W+w0o4
RAha3q+SbmK4mGXdPoUBYfTH9DDvqilvUAqcFFNLo5Sln10HoIORwR3IzKZyG98LtK+oH/kRIZtT
qO8wvagXhHDAUqGUyLpQtKIhIBYxJTTqTJ+SPHQbHaG0mNeMN1F8w5fSSVhCcifFZUAKhJt3GQmt
gHuipkE6tpeM4xZ6Sy8Psq2PG6EBSyEgzVd44/T6QMRmopr50bldiKb98iRbHhnIZPC+fJ6xaTkV
QP2xUmrY8DjLjz5YToOQz8u4U0+onJmirOzwDB2E616so1sG0svyyCHbmdvYOaNIfzDfUcn84Qxy
EpD7y41aoqTTDWYNYfkMon4/uAaxSUcLJJ2fFgIcvQgYnc9aH0r53aOcFiAPE6wqi/9yS11Twmi0
WVkpizHAU6OaPeZax+IVMpPvGR7t6fwi99+HdeqSQOTYA6gSovWimf9wvB4jkQeTh1Br5szUoqFC
fY04Bj/ydhHqhlmb7xow+O7ZZhN4VPCnJnQTNHOLeQPh48CBKvcuv8eVf3ENRya27qAF9isGwmc6
d/FgAUzTWS8EP7ql08ap0vneeTc0tsfzqqhGc+3QAI09dDhT/P8dNsh02mnAo8mOnE9N1WUwokpV
ovMlAcHl8mFqfd7/Je82U5nenSZB5tCKIJtoICqotZMVEuAWd3/SMNWBAzBGjwTdj54ushJNP7Hd
DgsAqmdra+imBvb6d+mH3E1LxKg2nuM/LR0uqzIa7van/AIOUJ+cbz3/r5NEBiepaUXa6yyFRkTp
2ykHQr37mN0YY/Qw1XP3ADfAl2XWlxN0gsrdhRB6A2LFBM09cpL+tgpOsozr6WW/P9g4pK4VUzOp
zjt6EN1lD8ctcIrXRC4vwG9XULzBR+309c0BF2cqRJWgU3+LiP3gvZZAtUW/QvCenTo+wPHbpfM2
TrlrC8HJKvV4MO3mYb7ghFrUSZrLCwLRp8MmpacG6deENt2FdAhbgwBvA0JM+3SqfbPjGqsj4x91
Hagw9HKiv8fTakru+UyuvVMpOEyJ7aGL0Mohu5VKoomgka9gJv1bapzkKD8xtwddoXcS8V93f1b1
pfqtpEUGclzveh87VW4kcj/p4Ouu97v/Kya7wT/2nAn2KlOsCtLmApAxucb+yzF/SFnKGc2Y11uu
1XwC0/7EkS7yBoLsvREyK5UuzF4vpGv6R5AqRmfreWL6MVqcdSoh9Om5YU6scehzGneVuJZM7dmk
caE2pHDP43+CI3Lh8Sh/0L/McdkWPSjU0XspdiWlqZShG2iFgevqYJ8flXUz4A6x/72elJ5NgdpK
rNwq+6rf2Jer+Dlwij2H6GPWAkzWS5hT20/HzpThUNyusK058f+7tQaYyBy+N/IZuabh8XeQ6wXz
odwfL89ED2WaGVPJcS0A+4FoKcuZkhamkOHvBNt3r1re5n2BjvI/jI2Ku465R4jLB3O/GXZR+dzb
b84ADpL15VfUjl674l9nI6VOuR0dXnOvm93K/9XzQmhCN7ktwK9esqOSchczmUpHqoOZkKJdy/Eo
UYItaUXY/sFsW1/5H1LKdEsTsE03juGooHQxa5F6YICLCid2NfM3FkGuNoGSCEEusrnBEwWyhHX4
Iaa2YQzC8AKTBAaPXzsCFrTy1FNMSFd/TUSB7RrIwLLhfFsFeDb/0jXMSas2QoV4QJ2fom4M47mj
6cvP9eRZ7yCGJxGajY3sVaH/OEs9ESG6Qbs1euet+5Rh1R4D57YSk4oi2m8eKdmZ07H161b5WCcN
tsd6Kl/fMBNpFogHzeyCwQZhG9CiCUG/dBFZhZrn/07jziWp3yTU+njSb3Uu86Ic1d+0yvZxEGGy
MzqIlIsS8rJKkNIrLupSQwUDRTR2RCIeur+Z279FARqMyglrPho4gTCJF48N1WZTGF0qWtOQFPzm
j2SlWq+FZeIi20FvhYY9B43NUbaGR6ZkS+q91bnpejUJqWITfS7hiMYxs2riGnOtM2Xwu9IRetZh
vufeDkQCeNYxymi5dIRuXrdGoVAuf0yCIcKdETlaknc0VirCxJAuoE6XNVfbinlqGfmdKojNTBI8
IAagZt8lTv1Xn+PlhzxyfycaZAhq5bEGSigY9RKA7Zh761vdHu6N29AbOjl0W8EibhQQNo3xedpD
th07LxG60oAouOSfyuYOTFErYDRYRxuLpcbC0g4WkhCdh4IBAoHhWJyBbuk9Lq0kM0qEQ6YNxyNL
9C2KKN7HQZlPC0tuOOgoVT4V/Y/bZVBc1C26VAdt1BBH54Eb2m1cs43fsnD5SzEse6DXRzwEkNLj
ODyoFAMtU/lCkHlklAoPmoc6NhnvDNemlqO29BIG90nD+gpSjv1kh6ZF4XzgZ4Ta73flNaogrKVJ
q13z2m8X8YIB5qivgppYODn7PTyHYcr3sMIPu7QbBMDZ5q8EegMRCMXAaXhp00iKZFo3Ya3fV3Ed
c6PwMEWAxYgofhSwjSCsPccy9VEOuztxPS7pKR0I4Ya1D05EtNg2B6pvCRuDj5eJZXfuoHA7Uj6J
fAIs7K/cvX1NNJANajrl9AQizqi+zfVGr1KsjdgbDQACnlUnqwyUnH3/4zOE1Q/4Gbteesus49Oc
WUYn85/4g4PzgtxhOXZDA1SWj6eFQnlK8cxPPvcrg7b8pYZUjmcaxLDj7URfuujqSExjmg9IQjDl
wt4/7oBoGOl9dawb55XFfQtu84ggK9uFfHqzqvmowkBx6CG8QzZ+JWl+gPHzAVQvNvaXboD6KXxz
lh5QaBxwXUQe9PhmuzF+xvNYrMXnCPrW6uenYfhTP8OQmqay77yK/v4nPYmertpzcWlN5bKcUcc6
RfJxGwqQ3ynaF2uUoWdSTo0IiUGxamzfmtZcuPbavD7ehY5Lr4AEWAmDuSZtlx8Ro6p2/E2xqusL
T6YGv+SRK93uf8V1jDVWKhb1BHn1FhiZx/ppabDt0bcnKgElDF3TYKl5/aDop3goB0rqML4d0Qy0
69tsZVB87WBscoyKernqKKPGsIO9htxmM3eGsfi/zD8XWfpkzfpDioM8LIkOfTLXBys5Ser4n82o
lK6Pa4UYtOGj2IpwjF2dul8vFxbWhtxkF2DlBleNKOdv5cfwFDX+emFK8I9yZkpfI7xQ5B46IFxy
TE8KJnYa/txOnq2/eyYAky9lrpOonBD9firaxXbWZdxsonK4ZpUlaTUtnSg6OWJYidf4j8lOEiDC
EXvxg541TMAmOUjBdJX8UVzLOz97RRLtJbkIxqAtw5yQKrtgjOgbp5LnuZQKhzkKGnHcrZNTgIJE
EXUWuaW5/Db/J387D8U4H2H5/0/6tyFMhk8kqK3t20pFmSIKc+iljBObEWHM+D9o4ASGywxA4m4e
6ZiQfTQ5K8Y3oz0EYC7lKgTA8Y1ffhwrLLASzogJfnkzpZB8THk7/hMqJsJv+mS7Aqw/5PG6/X1a
F2kOlF7wEMIVbtkap71YF88iv4XDRXFBsChZlFQsSIoUwag6PjbJmoL7nQdmfLPg3/WCz4RTLe1/
1QB9V79/yP4Pmx5WkxMnKlTyZfNCQektTJbMphN43ICf2TAQw0opRjQvFL9aY9r77xA9IP7exZLY
oLVIcycv5rdoK9tU2Zj9ZVG/fJ0pOyu1E6KsSQVSigfh0w8lUNCQIFuj2hxX0M8h+MJS9rsz5sip
RUDVn23X6aDR1bLYPFvNncTWvjOD1vKDIAC6z7HBxRD3bY+VDtFfO0auzTvKOBhyO3CYH6NZ7x0M
pHPOPAupP1NnwGA3QTqMA8IjY3ewrFJQNuza/Q9zA/Z8W90oKVLDXc4hQV2y6nsl2GFhb7JyVFbx
Ecl4/rqVqIc5IQh1LXvNpWVBinGYuBY2+qCB5l7xUsmjMbLvyA03tan7HxvZoDmOeqA5+NvVadxn
+10ubnfdPRbLx58mPrJ3dvfUsHjYOYaV/s0SKsQGwtvx0c9XahlcuKWjJ/lF2W6AT6N5jc100jtr
mqNKLCa41QUkDgsaxtt8EETwg8OKEHE5okYOnqUTrXULMBS8XPOEadaBPwtSSVdByyoZKxayHVaD
KNb5D0YXRIyev3lhQQEilrLTomWcHb+QggyfIdqtFgODgElynQxOUPCBMo+sKse4Prt8T4SLAFhO
MWkzcUAXkk5uM2MPEgAqfek72hoiuClw+xmIcDYIenSXsnObuDO7xLNFXRjf2QqqIRENAC4k5Mvj
S2EhTJEAwaiFZffA/+wNBgLoUDJsmCEUZlnXcfXFyTv9Js0RcHjiSahSQUZGPoR0W5bdCbMPIIWJ
lziBRR3AzecZ1ReQoC0U3bHRaVC60R/ZkKBuk5Mwp5I1plmf2l4+SCca9Bnvk9aPmjPBg7EhamJB
Wd40dPJaDrTklTaE46+4h3lrsbxJ3dFh1GnljWpo2AILkhdWQSBqN6L9kzG/jwzBc7/36i+3hL9y
I8SF9GvNrvGmQSdP4dw7UHI7n3rcp9szXhH7E+2RKRcCUha7mOnmbg9WO2wCSkvQaNP1JfPJvfc/
iEMWYq/B3mLN+9lMNEjWcoF439r24lxgh5rEWWOwKIg0+r5WhtcKlzso4T9vT7s9fUDxdLu0efHJ
CrhuI5kheDax8fv9Wz2Xp0ahsl5eYOC+VszVmt6QhAd6Yvut2avI9aTlH1RPoIXUKhN+pp5VEHjm
/51ZNh2xJrxgJYKpLXpzZprQJUH+OVR590iNZpyLtodE3vSR1yh9PVGH4bTSuo4OqCLOqXCP9jTE
xwxyO8VqomqbFhr4e+fdyI4Zo8K7oYjHqc+ZZnLOWYbtZiPgJVHwNinQ7ZQPH0gc8lW47V6Ro1lH
vQ43puYohME1v0M7h8z0tpQyo+VmJ8creWNTpxgRsmUXFfd4Wqx2fwEgvbMi1FkK6OF7oQ3bY4XB
EOqSSX3Ym1IpYpYfB0GkbQ5ay3SFRiVx2M3PV+OhOkWe3CmVVUueAQKZgepuAWRRaM9+Gf+Euuuh
bhIz1cKuKDy95/rfRiJ19g7cHUtKtLfLtQK3q4KgoyVQXEmqHgsooH0Pcsfd5fKSBJ5XXOnEeiSE
IKHFyvccKNbX6Ovs+/kKzkRof4AEBqMIU2rbGYc1fVPEUcWgob27qxoZXqWBlXms52j7rwPzt4FS
mSUGbO6t3szFNdTJ0odIo/FiWwfvOk4m8LuB4pUsL42pHeACaLZh/3yawvBqt8sHCj80RNgnq4R8
K2ykj17aUhjWahjflARidyLljZqDUtHjKTJUKwNjrXWoJdCxDsKSAlCYyfth9a22hiRPUYNEfcqj
HTd+xZSSFbRgJSqBu5toKvZxfTo+w5Dn+usKkWIraq+g85cRiUgKbP2BzOD7k1D3AxNjuNcvSEVa
+bheXtQfrH62VOVIuoncG+Q9w5Ws7BgRBIckqPCbbupneSMygA7YOejIq9dgiOhiU/pporATB0Xg
SMYbKYI5y67FrCwGV5iP0Kxibcpo4aK+8GucLUZmXW2re07OP/cN/nBQyN/4j5PKtn+hPMCBymx0
qyf69ZdmuJmoWJ8fBDltv9se1QaH44CdISWtEM4PLTCSF7yEFC8QjRZEgFwZZxK379sKtqcGVpoQ
9zhTFzt3A+bQcMi9tDIEwM6VCSqlUnZZAg79LmpGtdAqAzmTs0OeNvEcq1+genzVjJRZEwt6Oumz
1qg3ugO9VZqvEhkjXUEZGIYkyIkojdp0k2y8inmPe/5ACn8MHNgwO2CvV1Sb994bl3EiecDteCVy
JJdpnf8FZJzuFaoIZX8olMmvotaWRiGYg2x2fCuk865ToBJ6u/jUzKDWUMi+1vuA/ICY3FfY6Eci
TNI73hBR5NqSYFGK6+34iYoFQGB2TiKmyxkpwB0yWGGXn4nvNtTrDApRG2xrz/SgxIybkozaSloZ
UKQ5PT/KdmA0oGdeyO1XLwLHCbp8g7/oOpqxHqAh3yrgWAx+zSfkg+ulA3yOmDm2ZY5AAoqOTXRf
xxSnwVmUGhxHCNHhJ/ly9iuHtFa0xAhcN0dX0U3AOHvwH3UIOq42qWd+anGzWdt9cxnaNSuaSrqs
64bDP//Sm0kU6tUuVb8VIrdyCifakrKsII5PCxNFT/hYDWwITE+S2SkBiP+jUk0QQHzVaci4frW1
tisn/sUsBSFXGY1wkESMwBr1/ftuyplfCXaOV7ETRkajmI7aOwIc91hZP9FdGZeXZ4mnfXYuJy72
TFfwWNrxteb3BzEY4Ps6GYDpZ6A6fMTlUsdPGlzix7oNbiGEzvxsxcNinN65ysaEV2+kVjSN95Pj
ie2YnzIwK0FfG7yu2/eY8f1sCVBW5TxtXqgYSag0IyCOiIhZqemRDCVBBU57c6oTYLgxLW9HQfFg
1/UgNy28ni+0ME6KknbGD4Hjopao0+jqQJ6QRsh+xTyQTBmTQo+xmIsyHDr0FAZ+ctOQgN552IeY
qcsbWsGe6ZkoyAHhcW5MwAUxLSKEOVc+h87WVAhORkDx1A6Cep3r7B9KjdoAd8O8/SqmBGkmaCn1
DTmnG+e2IbVI9j/NXnOsRCojwrBtXhutv0zck1aWtJcbU7GuC8YC9RXu6Z17V4nPL88RNGxBi6RV
1Kp+SHYoPV33zEFnvsgnrH/80ROTMV7ssnMmYI7dGQnd9UCc/UzRXiPEUBeb3PjTDbHkjA9stNma
eEAp/rTnpMAiOfVXQkGmV48zli92VCdVP89ECRBfepPxDmGr4gP6J5UKh60zLIPQs4K+debk7oJx
eLpMzTNfOJYnq+i9g6OLFiTvfgomTfgmFuIgJKbp6YUHyygoo8Vh2/B78kzPj69uMEiC6c05fJYi
vEV5JD79phlUKsyGlFyxwTzgbulamq/HaHHGLYeDHN/8Rw85PzfOomD06nRGDzPXXrIXNrATeK0m
qAqplluh/rK6qx7eoofBeErDrMGECDgggRercPdKAa9Ign/yHQHpIo2zB91boDtvSy2Y+obBmGHK
xEuzA0JjxTQAQ5gqYEVSnAVNMofIr3QtnmCI4zpWJSDDztVFP0qNnFO+6Wzmu9DVUGlJjgrcrPe4
25TEQbKviemAATQuLbMy5ThsgSaqg+4fEmbD+ECS524XvlL2X5RYwJnXSez/BjJ3cv5wJb0wlyZs
joMGLhSewOqLZG3+Ume8kdIvvV1ppifmVm1/b5MP6FtFbYdZYZY08JomNfjHxMgaGgfsdZ6iH3Rq
o4+ZeoIZxD2OZWRXvceHr5VKQzYwgTdDNsQKuq8BChl3JAdL26mTrjHMQ6f1wD430hYePa/mOgxq
QUbWQwes4du1bgonSy233E+Kmn/+d8MWxZObHK/SS08g2tA1U2SQmEVpJh7TuJ6UfP4stPDBKdvB
rR9WqSOLv3cpOknYoqR+MmHSM8qi3gC1Tf0ADvPB/IaElcCXQCNDcmgiYRCmxn2AQbQPyTH/xNJx
k0lzzB5j39M09rrnKDYFrGU197FjYxZXzsim6UHsyXoL+3lhSeR8tjcPMmBKbNibYnIsyNZa16bV
uJ40tgJwb/0O2x3A2ojF8WEq1+Qh8l3zNj94WJGD0WbKx0hWTdekHXAN+8T0nSSDDV9kKmeOCDM2
jPm/XwsilD/KYG9Qgl0ZuE9kT6y6CUrSX0e988LDsaU/HH5ROk19cCsWMo7DgLEKsbg7am/wuN7P
uYHsv4WPTl7bTBrV945QbuEw/h/Vbf9ttw7hymque/q7K+a1l8tWVQWWnSA+C3/NB/431RW68BJT
ALwsiPJvEd+QIS+TLzH3F9rwrRcPYJxaMk/kRw8Lrfur6zEgPmt+FIwqOsolyRvYKAcd/eNmDtBL
IbzirlxE7pCYa8S5VlED97QrlXTvLOhjKw06+zbywM12OD0+Yo/u89W/ddQPd47Q0RlUQ7FSjTIj
jr5JtA5jid+kYhpnHaSO8hRHko+YLZ1lQn/NxXPSTfu5YcyBtYTBt+w0kTCSq/qD3WPYE9gHF5Ea
8ki5EYKHP+v9CN204whN+Wivdr53gwenJfZIkFIyts/2X9rmZFmDnhOoG8L1pNMvmIOmfxBcTPdI
BZhfsn7i47tnDq3ySB58DCL6Odt1m+of5cUvZQG4B7AdUx8xWWuy9k6vnxxj+PF6Ef0YXuPD+iW3
wQDL6OZtE96cHP7rik0e33dHqivdbENYzvqIHPn0oOWsLMLcQuokYvFpclNF4T6oxiiaPGEURj6W
CqI7B7JGvCv5V1G14ppOKJmcVzbfiDD3bi1rPcqEE8Zq6ys720lbK/pr7IJBI9C4hl1Piontl4bH
tUbHHk/epbEPLWVULIgUelmWEJm3GTQu72H+kj4ChBmvU39gJjQOyAgCg62kz6xXiicfh/aNJS6s
znIwebFyKVPNI6YsxJZZR5yy+feFQVZ1zHzV68q8KfSeTRDAUHRfuA5Zno0p1yRAIMejlz2CUd+x
2JjVNJlTm2BDS7MmyvdcCpiiYgTQLLImVbR6EwXOg493lJXUGDt3TLClANIIwaeL/fTCoZcaWUH/
61IoL9pfW2+Mp/jVn0xwPYn+rDeS0lZwVi4PxRpuX2m5582oLv2GfgmdgHdRJYfeGa+7BuHa5NkZ
ZJ3l1gROu908f8B0jw4ur54C2RDZdI26/yU9ggD/nZo1YLjq10CmMRAWC/4mQtM9B/oQXxOOeLav
o5Hvq301if0xhEaGEgsPTmr0nmue0/YMWVFOnZcsuoXEZZEMOvbGUIy9GMCN/3lxqxpyZ25tEzjl
90oF6M6uiPopDe8a+aY7OaoqF9xhdVk9eztVq8YJzRp/ZG1x2166HMkp1zMkRCVv6K3R5S9D7/8s
AKGKbyPPMRrSBWb1o9bNzlXHo2m2OLEmrS4sAkI4FEU3J1knsKT+i5Vnqnmli4xfNW++zE+lfQyQ
A9hw1cMLchYf6IUU+stj5EAvifv+HSRjnmxWi9GTERtzxEB7ktHHZHAQed2q/Q7/MM++PpVqUcVC
lP2C/s03cWAg3Sb9C5BD5oWDcaT5sWK1vmHo51OTwtA9LIcCJTdSdEgbdrzzCx/ydUGOkEDM2X/t
fZV9su5JFtMYGjjCHc+SxvjcPzi3U1tdiuNszXYRgg6V9txk6NsR8ihdb909Gr/WDhyHeCUt4ahn
uzBU5sdTIl4DvmEHqb35dBsHpw+f/VAtxMWgxLW/LgHVVOjid7ANmWf+96QLTnJLaIyl+Pl+jQLK
YRmiQq0VGvsn1Ih2VajDo6kJMZZ59gmaNcFSMwbzljcjkH/Fb2RE3ozOx+jr7EcfTPsfRIj8EBHY
Ck60N9HJSU30JiZHDxSqDGT5kH0BZCraDNmCNquQBf0QmxkR/zdxSt4UoxqbCYeurTyQTIPIOKa7
sgWQjnhgf2hXNuba9/Nlu2ZQhr2gazSESBNalojL0wb9vI4afbPstpvmlKv8/6t3hB8TT8gwK2HA
NpHxglZqO87HRHbn0NB2GELBv8McdpaZb8YDyTzKtPC8bs5D0H8vJbGq6u1tHt42eJg7S3tfHmh+
ZonNyyZURAnLYqg2ftzRl8yvx8kX3xrzSwlJmIoFlfFGSj4CsqXljOdUiuh6lfUZnon/rNFQzjfR
ReUdmaQXfwSsN8HdcmDaPaREYE+MQnxJId1fSt/fFKLV/jclgefGNjei+yyPrIwJPY5j2nWTStOF
5vc5SuBkshCGCR6Uigbn35YzPArgaQ4Sr6xvcu7CIrInAa7HpSnme9uAwbygvi+mpnbjZZ0ShH53
HE6EyxZXiUnoOwgIH3yDyTuNgPmKSRL/HmzxkdAkSpPW35K/So7bCwH5Fr2IelLECgEiT52qrtjA
RIRQnkCAMD+1QXTf96+POjX9r69pc24RTX0uow9iVtS8Pwe5WaU9V5mzOSM2fvFXfDLQHA4Hqs18
JlwTv0h88Q2DuMTeKpNpdjB33Pc74cmYpnUsxRmTu+jbY+f5zNQHUzH6j9GpzaLC8+8XUW6XXb0f
hmP2jJH9vitsTIffZsAdtGJ+yLDYGKmoEdiwN6sm0fhpKMdsHanfCZW7ALSZvoc/BJge+7Vx74vU
lNQ6PoMmHU8s7AfIRjKYb2fmX9w1DV8E0AtyCeY1YSwdWv/e9e3mSHDlpDjveQ9cRzuD3HfhUjPo
1RxPdGpDZIyv2wXeixhR8FD+97ZuTSrATATS59eSEXXnueDOiH6z5RgjFs/oPRgCTCEDQjTb+D2e
Le0SjppZNBaEg4q6c07Mn8xsDv/dPWAXBEK9TZtaY4LijMkWcJJZ+/Tba/9Vvbaww0pkESmjPKvP
FsZOD3ZW+DFq+ckTX4NukCWwHvz1xo9h0DDBVoSHWWOa9j9iS7KN6NguN8AESmSIHGzOiZAxk7Zs
4Xc7VytZu4sStrg8JyCuEu8lPkNYtiLg4rWfreFXZXKBwCPjEHEwKmeeRiivaAifdgs65QBbh/M0
uryb2kVszBidTRU0qn1reLo1zAt+QbOOosE4QlO3Oag/PogZ3XRCnYX0nttPKott7XmTDubpvBQx
uOV1qekgh4B1MkTaScS7nJigH1jUJGAn/ZzWFUcFPsty7o34OUNbGsvLZBsJMD3aKYkEKayanvqb
SMsEXhslkKPO5zxVsLXSrydT6rL9IQTuQQp2Etzfp3qpJ3oq8AjCKadmPvzNz07VO/87kTmc4b5h
Hux6yhTMpVRSmzPvivYo2Iec8ZKXLo0HD9+JrDNSkCqJ4X0onedRHDgYGEcSln8PO92BT6HlNkPC
EhrfCZ1DgIjueufI3ynuO1q9tMxiXNk3Lks1NfQPHMUwfirGDpuctTy03sYMdYG8vvAttrRUt57W
aQWiSnp7//pOe/sDcIl+rkA4iQnCnR8tasuXdJry00WuucJdPMTavNhba41CHNaS8FCP3bjDkCVe
1wLOUpJrKKWmeiy2WHhBJNr8kplDGC5NmQrmolRofA0GNmKeJZGeMMa+Mhy3+5KJEfaBNvqG7o+4
kS9V+Y8P4fPFpt5Hq5WGJm3j2U89eKW7i/KA9r1OkqvrkUvVz94ZffDnjV087wFwl0ZMox4NTq3K
V8sm5trPsiy/MAvB27GsqIfnIk2vD1aCY2B14UGcsZEGJOzBq4XPM5wswA/pJlYJTdrsdOm6QQ/T
llVdIsK2IU3NwIf31Un2tz7kGKGoc9uVu69dqMLLG8Lpk8Q+kyOIQ5xurpRXG20yuiYvNIpbb8Ic
+dY2G9qp6weDZh/UO3cNQFXc0qrPV86+U1TqOMuMy3KJmVpWMIwz/GMxojZX0WFGoRVd5IIRnaua
XSFLH4x7/L0OsCTUa/onW65T0iW8UNRdj+uPviNAGEtYPG0/DArZ8bLmnMWlcqBoqHzsAo++9pkR
c5WSlSQquIEhfJ4P7ctwauDv9Sv7uslv7Swq5rftByD/acSHR/Pt+6ZQHCPjMVODgtP9ztKbTtZ4
1OiqiWqQIUbpzYB4vn91bfjuZqwzGrR3CTYWBGwjjQWUsMRoNBKxjs/Zl0JZQUidE3LssKD6Z5lX
CnCp5dfx57F7PwcZo1LXS+MyYO2Qj6DfRy3z7DJxXWmQLjzJAZgOdmtz+9lD3WDN/Yt5Kd//PDQg
LpGpr6/wJpJSc/NQPCbTt2QjdI5pNRcZKKtYYBhnrdzyY/+/EQh0dtMY76Sml00r7A+/aNhy34Td
PpBlI7kYr09rbyQyt4O0OWpAnV8QEcv84zqwfqLFN1QPWwo8lGntMMUu+HPVWLP1pZqK55U0KXv7
IXpQQdLIISss2jFvbiUpkOu/QCMFYckQDI6OfmBiMAo1lHWisrJu5x+RIgUTetiev2VHf/GPPkXw
TUQVN0nsuUzrFAbOCjaMPhSV4l7AN2GdbPW/Bpwp+H6c94Hx5Zlhu9b+4tLZR759CEzvAeLItlUm
WSe4tgo0JPn4EC9CvxIgkzz9vjn5DVMQHAuH7O3+4qmu8sd7oyvHB/uWVRt5Rp/9tX7D5s7gbrz1
vFkeBcE5qM/1ZPcFN8DfW6vCvSO5+1jCuJDVNgeNzPmq3w1RIZ2lVoT2Dlrtf4WCjMdKz0uh3HuF
11Y53H8vI5rCfkmg034ZIsrARNOHjJhv97ctndB4JTpK5Hh4cknEuNBPqauw61rrg5Q3dbka6CTF
IbuIxIWeTdQiciD+kV/N5jRRI/X/zvaK1dBLmqaKhHX7TZXtW62kQEvRYDCO3NEQXgAHJ7zF0T/I
o+qIoHneSydNrNoYQqcZT0cgUZeQ+QyP84TGOIAR9puc6MEBYQQGuWdLfP1rzS5VV4r+G8e5KGOp
8Tc87KaS4lNb2fm4v0zvZM4PbTFNMeY//RmoDxLFy9+JsGHK4TpMtKEvDeiFI5TFrm9lx0agzznu
2j1F5WswM1Q+PSAeSkFZGug32zuyni+hkJsNnuu+pDADJifET52cQ+aepe6aBRelEkHanoo8hETh
KXy9uIQV0cXM3NxUKLhElSoF9KdgKx/CGfUMON2m2YLYnWccGtPNjeZ4m2ISsvAaVSnhVeAhM6Rs
JhpkDjSkbqqjA2ukU8rQbpVJKsvodSn9pkdg/wWi2PJYzl0+mAMOflLnxan2B2gqruEmq35BT+2G
dwPgg9Qh96nuE9p256Lo+c5zppsNJ1MPq/IoTa1ogqRF9ADz5LUpZGU1RKJTv88q/gWVuGSPSmaq
r6YCkXko6TikiqMIwLup/Was4dA9aKUHa0jFJYFdpsK/W5T1B4bRm7bkC/9Z9gUVtgsYHHb9ERi6
Lb3SQ90FkAzg5auqO/Lai1q8oAi0FsxvVNjJZ6IYG63+O5Fiv1xNLfEao/R8i37B92rjmUnW7m4d
B77WCUysTdRTcT5V7H8+VKl4njr6RpRB8y4srsVpTnA782WlLVrcQqvs6DWWE0ErD6QPYSX8eKGa
FkvSpPP5xmhrWCoD9ROb9/arzLdP5UQoqhFzotyRNsZQ0hP0V2j9fNqpzv/FvCfaSEHhzGF6L7ZA
hI6MOAEihKG0OGjCV4sydGOpO8yQSqmFo57A5IKoDpyx6y1QTPxnLkwiaClpK4fAav0nH+DG9Szd
5jicxnh7e51XvHquvvIjwzQ0mvj0u8lA/g5kEi0t04fjgvTJiLxeWXYmDDAz/sMcjLeafG7qijnx
v+8OazzwXgUWq1A8dhwePgKOOgcfU2U9rv3iGhvzYIC+xTipeCN/QQ6HfjYFkf3NeYV+jCi8Ok9K
R15EklxJORLsAPFMP+GpnojBDP5bvo3KQaF9rH+ab3botYRh8cDY710t8uOU/8vFP82QUVgE5tyd
PG0WiTGm4IM13AaIlULrLHTh837fAZ3aahGOfI1BwY5D/ghMskn+RvcglcbzilWZOQipLMuEg09q
Q/BEggHMel9Cz4pdDuP286hXwuDqCN44ZsUvCYR39YWn3zmZ/+EPh91urMGly6UHTMVVDJJqy+bV
+ckrZdrWEIEa4Mn1ygIxeuu05Dq9wq5h8gUhTTpR4GVmNO7/eor8rVrKLPhCysTodShNej2ojNLU
8rJ7yFNRlGzLyDSL1DthcrAPtL3HdyFwYyaoIW/KutbZ2MJgSEgOLQ8+cKT9uXjMIH4QH0FJiNPh
v1d4j3WPZD8g5WTpmSZTmbbpPwZF1EUU9eLxIicbILZQL16WhjcnKqK+SIUZI4SbkC6Li2nzjbJk
VbPqTDZ9Ydw+ochg9kYL/uDFtllsHb/pB6TvFoQh2IQ3Hvc/ckc6cx/arl7H/vVd93xrpruip/YP
1siZhWNyS2CZJUjfpglpROaxZ6HyFVW9ILCzIWh+m8wPfm7LdGdChD0zJ/BLv5kGjWPhIyaoyX/u
0ESAJx2pIcgwnLYpH5lrDrkMkwWSM4KK+zofNfLa1siU0YeKXDRd3g6iTONeGzmwzntPtiTdV3qp
WpZeSDPviC0SOunDZ4bwXyKx+oXEzayEhW+3kh+r9C12nNJoSE4EHIpbcgkPqojzw8kvjZBXLjNw
jorybuHNWXVxhx+x84UORYHsz1oNu8Mpi7gbwosWfYFbpS0zHdQ1bM9a1id+CuFe3wshhtxqd39p
pIZ3IvK5Xzml0WCzenUSTgTJXMag5KtjY2TqxA7j3zMBXP9LQwKuk1I2KW3fFDbvHQFGvBx8yNMA
aQBRFRy8du3Vt1xg8urlWgtR0YCjUb/kEPpP3Su8czNHFgOx3qVS1pp0A/ItYPSfXhFG7bsIHbHM
uV4+kyCjqDsjrKAPrUYun4t+jSJMve8ilRSVR/xN+Fnm4QSs7VUNU+ajfQTNJiKLCSkAK3XkBP9A
0Kvl4kYfYdz8NHrJPpt9yOmOoRlfk5YiwsO7TIHpraNaQiYJMFAlnY9OcdpP8fybyTj35h7CzV9a
qSMaABW+1YElpeOne+FvdL3Yuss73GaP/IzLO9pgtmeCS2E8tPmNJScsJFg0/QJWddF7HIR7hY0G
NDHUx5yiwT6qsDGqRbMrQB17cxtzXN/iKWgq3j3xBiMfInRKM1X9UAgV6/3epvBoUWkw+VEZBqas
KNSfVPw1PagjsPHQWFF7TE6gi5j6CKm0l5iqzSCAG2GHR78TFD4nZI4LwHYMMyUp4th4ww/TPzis
dB+BpFeJtbni8cGY4HkCd6gs1S7Ur7Y5EJemgrrD7knfJIpilTsYcOYJ5LuqyDti/VsbseCwsx/N
6EE/m3Vf2+rdJjf4gQpfDFyGPNaHFllQ0QKaILdJAikqNOcRrkarBiVjnCsnqydpMqlHdj90bCV9
3QV6kKyVsOZ949iLSmJIC8jSUNU6ZwWwa9Mgt8XI9a3rot9Zf5LE2ZjR3wcjjImZU7KM3KU+MQUR
vKaLV7ZeXbZ9AaCeliQ09k82Nw88M1YiHyWvTsN5orDMoqo71doG0xjqaFud9UB8PGYgZrzWbzru
qUGs61fq8+aICTY4140sCKV64W5qerQ/UnD14uolg4/c+EuUJ9FP1L/7/Di/NPgp7MoSTgFr5cUz
f8kmOx1nVRW7YSN91S9tRH0J+nxHKJyUztzZ8KzZCog2soogVuvVfHMF1eRhq0DDxdQyRFDgh0ER
oWxRqD4ZjbglaWMcMlgpt8iM19z3jGuJzfLRfM251MHFiAIU5T++fqlmj/JCMySY4RGRW85ZdNeR
cUn7EqUu4iT128nE753yl3h01zJi6L3jGphpAxJQa7nFwIpz9TlUUKp/bglzeSUQwq99/XidLGmS
MWyXwFcc3WXQSPj4UTpJga+zJHoWWFmZS79oe47XGFS1OVGAkW9FVfWIhPjoEk2Gx3X+9F3OPfTU
wH1Mb/gD1M307zLdNSDfhJ0AUIFRvH3WlW6yK3KcFfr+AHKwsLdeE316xxaW41aeVH1s0mAsfFBd
b0w2RLRViFY2YWunbTeHN1/N0+U6O7mTgDeZdES1aen/Ot9D2mnnCx8BV/c2eqdCw72sgncEk0P+
dB39zHhCftI0iqGrC3AkQ2eIT3WlxqlzYT3vDxKeMtKhXkT6e0npmvN5hf7Wwv0fy/9AEPf+h8B9
z54M51kwxd3EzINWeskGMSxYNQOKIqjLBEH6nt70Gq50zc2WOh0/L2H7sDxaGT3NcLcpbnp1Swdd
AYlhhogOdPCfRIjyRgkNw+7+HfRi2tB2cLit61RVw2XPeoRTdXZ5IWJMSZ5vT95b01pu1bPhkJQO
2L/tpMyCVQL2mm/gdBKphd0tyiwQLuFGJ2aaMj8UJYa+0JuBBVy8dQfZq2BLtLnWMGDukKjzJtp1
BvtsVORwYQRwoojIBUL7OvmWuCY8aJN8t+8yck7BHlzoZXpDAYYRGE59bcBy2AQaCORZKiqe2Dg3
gnYoAcd8N5l5/26RievFfbq46Gvo6UZhZsFLeZWOC+vWlTDsFKIpJdQedgIdl8Vp+HE4zKoSd/kx
gQU0VJXxJlQq39TPKqQzUmQECnjBoSVOn42WfXqlFNBTdnYXDBQam4EJsqb3NcCI/rwHMeIC0vwQ
RqRMpuVnNJLdO53kZeAZsN3BXlDHd24B6b6RyNBGvvAf5ByrB7ZEWCj4+F8tJFe/9GoLCAZCGGMc
tlvfelScDfLE4H+HAGrNvcVf7gf6uiKRURRC50aLUFeUtOQ1dpOQVZaVYfanR4SAl8b/Lcb/PhhS
2Q+ZuTjFMMK3QsFN4dvT1wgUdEx+DI6out3br4qn04jqMb2M7ybEz7MyQl28evM1Vpw+dXs9hC24
OHv/9JQF5WW7C+uzvP1YvkAFcApjll1EIj482xvzd9Lv9Yd4UyMobVX0b2XwKaYGhIWFb0ohzcas
IlIbke+JEzx8MEPbGDrtxMqu5MnOJHrdPr9/FbKc9H2M3fgGL/znzCzGsuBpEeTGoEo0YbBwdCFR
eX1Mm2iBF0m1anQSnmEouaSmQ4u9XGVHYLK4D1ANUIxrhpz64+cVa4x9M9e+G2uK32VhJWgbZEDs
gpghMAR7bKN0haEUA7OAK+SWUEBW2X5xHikQD1VlOgUEpFsQVZO1Y+TkkGm8AgyQd+EtdlVmU2ci
av0mAODdyGXVBd9wwqXXHFPO76Yc8rvRFf+y300g4xg87FCLHt8R9ICBlRDZ07wIpNLQDpDbCP4x
oSf/dmttvITFy75zZOdDip16v/IrkXWEGenBMw80mvCBVu/d7Vi8dK0JGHjn5hzbcsVR0toqRuVG
P29OXO9pYEcyIMk4dG3fbnx8GLnUe6xeLQJDYiW4zY8E6IUBh/NnxO/dOpbhUF2njmg3KJbE3XvR
Kv1xZtXnc42BAGDJ7I8FFiHOaex2u21JxgolJ80VDr8hYop1QMa+wu24o8BtDHAjpj2z/YXlRKWh
zNB619GYchVOta0IgKvwS2jppjfQqk0SSNfa/0MUI+NGdocCcgdSZFOUmufW8UL0Tje7CwS0UUGy
ATac6QAWVmcklqQFjq/PYRJUgHlP4v4uEWfV3+OQuT/PDikDN5aByWa+xUSnk6yuxCYuW2bFX/Tx
DIY95wsL4Kpo6HYJYi731tZjcXMJbxGVGWT008xrBl1VpYnYz+B0a1HATjAPJR1P0mPEReBfzE7a
8sBWUDHqdFUofnv839U1kR4gwsK/+0NntsTBwsHGeA6LSQkJ8HwSrqttpXNJgFhkfUIuKPggG5Eu
JFm0Iu6B2NV0WgV9PPBDx4BafAV9/SSHwAgOrW8hyVYo+oSHx6nrT3OgriSL50byJXa/Ry9YboGV
5IUdxbTW57nbJjSRBEqutgUGuoAD4I6XFW9eEOJyfuU1VBz5JbBDIdQHjhr2UIh/HgbmSNl0YUDO
V3Tzcc6soQEn3OZy+Q+ynAXh5Uppm1cpQYRIq8p/neL0HWebFRx48wlIJ6/Rm3bZOwhIhsIsf7F7
xuvhn+XkheIGtGESbWoifm1LY2aFzyt4uaLItDO/M8UkA0I9EYq2b7XFXj8cp1qL1KJ/U4pt9H6y
V1KsrfrP+Kv0ynFbjhneF/+7rEnavI/XfEA6c79vjazaox/kMVETNFE6OZP9CrYFR1WTkWuccK04
tC9VKPvgIrDMOurbZdKr7/nAT+EflUiGSyGulykPBlBPi8a7shGDdHmBHGE93TXGY30sxDgSEXdC
IEVRjgFg7E5qRZjxLZm6iZLNKxwL0vtRxooNSdN+5c2iF9BVg7xtFAmis20y6n7onlL/Xr0QiTv1
AxcK8SBdFu+uE5UidRBGXgsx2U21jy+OFHFVJD8XDFVYEzP2rjHCw9kW6f6LYukQ492b9LhzeVxF
5N5PeMzjGozq0HJt8YIGLyPNH8N3h17VyUyWT/+sLup31OjrSoCOhtST5TokaFhDha2Y8k3ehwV8
/HKohDlcW6ajRqH2hwE23Itm7Nh6PJDJwGoymQwlxS1Jb5RaVx1oCwWupV2iNhyoPEPUPgLkNL/y
INBtUL3mafMA7N7bijvzVcdMFA4+bHwPOzE/bmgy7xifgTT93ueXpeZcEFmVVX7sTOADxwsm4c76
Gp1GBsphWKiZD7WmJNKPAjt+CLBMs/UF4tS2z8/VcLz0yAiLA1SB6P7luegP0bF5d//uQR8WQRh2
9dE8Ygh6Mx9mbFSnc8fdIoHwcybkidBTmr+2wNEDyoLsJRKzNRkPSo+4/YYlOsHOw5pPdcUKXKl9
zTD3aE9ZBDAXKrIZbS89RxHY6tgkZ1KtLt4BvP1tD/7yxVfTQsUnV8u7kyyFxaUFucTG78D715dd
j7e0R75Ym+qfNtvuwYbK0yI3WdbK6PI8o8d5p4qOloWFgYRFoxL1SXZls+98tLeb1PDttaRTR7FC
V1BOEF7zsZkC/eqF2wkDoP6CdXnDV2YYI7FpjVaxAu1RktDn5xfTk8B3BPukhCwBScM0rTgFpEly
9SW4a3+f4MwEjwcw5NfDCmTOuXMp/qKiMHI7XbnnLddY/OAbg71V7ZhWke54/Gr5AAeY60C0KLdK
FtFgXv6wkybjbIUBBpMmD072MmKawXORtQARIDKA7ZCedpU1equBGvNCwJ6h0Isif2XiDswFT27C
DUZkyW2iUgzbz4jxYJ/tNNP2Qqn+39Zx8Uvd2wjT+QPrTcmmtncob5YhSHh8blqQecI9e4h4dZEy
MGo7HNVkNTlPcHTkiUbr62xD+78uDhX1j7A0u6gWZVtfWKXTj99CR0/nwzznePPI24bgFqTvnw+S
vY9Voi6+kBkOm1kj+KKmCQ9DvkpcqZTAE7uOEKnKALxRCd3Lvwh9HKPA6NSy+PmSgrUGVObl5BIo
arlAMHqUUNktk+KxcplN39Pjy5vmhwNgGWwB/GaaiOodz/n0PymY3xFTbPqR4P5v5loSK6G4a6cI
BJWbkHKV5wB0AX+nU+R4lZmptZk0dPzLNdttRsZT8R2XLTq/D4jKuJe6JsYnuPRvJUZBBrsoaFOO
QJc8wBUNdwU67VlmYaFz60xGvUxfG/s+eXywtz/B9kNx8+C2dalQezLIdgqZ/B0TRgzlEK3NyPAj
6TNwH1OrDFPz4SKRU4wIr0y2n6vhq5lA7cqEIYRNWGBx3wZ0YexNSSpxBwOwvQnU5eZS8jsxMBz4
BS88Kr5t7Dw0FmddJHpzTiDV6rcaOnQk2PF7/ybmCGKbj7CJikC4uilrLU/M1UcbJJQYv7JywNZY
D5QJXaM/69y1ZhzQ6ooEJOxeTlrIwG/wZ0DMu+TKXwDM7qElHYvVtrs+KLfytYpaSyHQpPr9U3uu
ZZkm4pqWzokvthMkvlOJeW89kWZCNIjbUCToIk61zfMnKkgT8LTPkKAZHrJVT3nT9BfiNaAoBvmZ
o+rgIzLal9KDhbjRDmq8jujvsbQ/O8KRBMbTFSaPadkGqjI4cWjT5pTRdDTwuRoBmpV2Yi1xF8b/
Ifu15sWID3ul68j5M+dJHrXcbC0MPDYDm5HfuvqLo5hB1KoguRInWSRvjhS+iYZXdsat2FTHOweJ
jn9txwkaBnfhWECHgjgteBYMl1c9WqIVS7X+CvYT4cpUVGNC6xcpJKjUrHYrhCBAedyojIAIMv3o
ElkYXOfq86wcqt8KAigKlnoLUfmPKZB+n9/vn4M3VoTzqp6PxAsMXqcGnb27h7LrG3LMSi9jnZ0O
MR6PeOAniihzxyWshYFnFKrUkdAhjPtS5YJUXskEFSqmNghGe7F+pc/IGuOWt/sM3UHXnoLSP1e1
cfL9RR27bB/QcAlDJijiJ+iwHE7LeJrgfMd4xmesPqceXhP0wo0jlD7WQu3NjGeNvLM+3Ad8tJ72
OZOarM1CgDG1HAmhXKCzIkAxXdbHwKGbmmhWdETfZQ2A0d2HamzARvVscCkbNYNVNfX+vT5A5qkV
vP8k5DXemick+wQ8zom1bb7evAV+T9c0SWc3rLyIvz4ri90OzpK3Eq0YK3rAn7ZvE6uaLiRkqu9I
qCZXHlc7rQKyTW8RiroMi3xmtI+aPhkjKczTBl4GCxL4rYd1FIF/yOhW+qC7+yLuSl3St4yxa0Hx
9QHxsclYg80Izc58ptDWkphM5LUiVnZW7A5t84wcK9kfCKJyvCEeWjZdRWlg9yHEQrVfq5c+ywxl
V7SX0cbsnHpxTALqe1KQ028BjUVALfe6PdTZJG92pUgcy0GqGe2x4vz72e9Xi5BwVWEa1Lvwt2TC
BKrIJCNbx5OaLyWan4iSxcQpz3MgWe5xfLMX5B7dh+rxUBKUogkwJjU9ZZ6B2eCaCtFeXKsemHhi
vRuFeIBw5omTYV2Pk7WM6YN6Yaj+mdHs/EniFv6KV8MdjFI7yFmyOnVOmEmmxXP844DJbGbW1zAY
BYAkjGjG9ygDruWtGIYDst16w7VrNatfto88YgeIxgoJ0Q4sJJ0JTi1ceEeE4KY2McztCIvZgyB1
D+A/M5+wzfCivYq9fZyjCtb9u+zcdUCbj48jvdIQOdnIV8N1Z2o7GnGos8PMRCRLpo/65Ul8tMhe
ae1Tu/HphVrDVjdHmuhndZtPFCdmMvXpSl0U1syY34yC0IWRyI3EHDy/eM46GwgxOc56+E+7MsUo
bDJd/Vgw1MiolxZFOdiZnJB+zG4xBDzSQtoAxezgcNtyb7AN+NEs6zPby/echZsboK8anYR12/VN
MOr649zBtg+xPB7YZD2zooTXE72yYjYSxX2ep0ZbUPkwBT3vV3EJ6bUJM6JsWYISvi35oIBj4Z9H
ITGryhhvHs5CQ9xb1Knv4EMr0Aoq/0XWm/QN9bB1KQn+PsgzINOxc9he4TJFRLseH1BHhwn9n52f
PDgY/CD1E8Syz6CtOZbzFQg6PHLJftp9v0xwSXge+L4BvBvbjDcVpaYoRWrleaw7ucBBWogIEnF7
/wxmdRkV7tsTWUYBg4lSUNmfAKOyd58pfgvtpd3UM5Wro9JX77z0y0uPpkQZGuL4sGNJ0Egm/xE4
B75DRYvtF+ptBQrugskoxlfoLzRuZaUxo85o9mSwXqZk+bz/gbSQaZK+DcO//yw9Jpu4kgHkpdtl
QIyf4VBh8Ew+pvEdmyEohmJHTuiJ7TC+Qyc2wfQmnTzriZTH3usBbSh+uLKVKgxo4ANIox/MfJd6
x9IwyT67ghfryRWzL/vHbvPW9XH/O5zQNg8jv7JQkm35S04qARlk780CBgQ6UYIGmRpzlQPVIdbL
EsrHtLa/h83k8WHLj2ftL48CAmGRe2R5TrN6BPWQ8W4hsboL17cUH4GeGNugslz/BwsNK92j74s7
8oQzb3rtcYi4sazQ0IIhlnW5lDFA52XMgUBp9QpWR2LjHTrn9Gh6q/3gU6gDyIHeFz86wYld+3RV
UJF20eWV2nyotYVozNdUSq9gOvQDB9BqzavrVNA3zBmH5KM2x5GIZfYaTCCO2G6S83bgjFXOByFQ
0pn6JrUxwUFZ3qu+9AW5xYY6SA/mNersa+Wo7Nr3edje5wNIQfN5bF/rREDMsmkiR2sLQ2kvKY6c
wsxdFeeLchMdatncqPlW8xfAr8T6gFw9V1IjW2znIIGZxR8SnCLKG37sy16/cBd0w4vQ7nFJwsel
hcqPAdpt6PrpwI+qH4Tg+EUamoUZiT+kmHYNn+DTyEoD7XW9xtyQvt81IR5w5hS/obOxRRWTTJ6q
tYyZ7o8nAEcjx+JJ2cRfNPxAvK9ciNKG5OmFUwgGutNgd3H1WnwHWV+G0oKjS0VF8N/hae+alIwn
MRVlXwyJTlvK7SQciidNQKtQV7JSJoDKwXlKo7GJxWym6Sn/+3NYEoeo0xOaPBElBq22CvfDWnyw
2tsFLHPgmqpU9K3gjnKZieRLCGxmKcQWxKckDeR+6vbimB20Oa0h/c1UNrbgBsj8dF2fHOXLt9CD
voVtOnqCxO8RGG3xm3MDykAn8tKsL+ZG574C++VogPvBRVU30w1U2cq68KD/NA1QPQC2OAZ8SXLT
/xTVWQ7Zh88kzjFhhl4JgjzLQt235YiIngudCBS1t0zgiRY2hXldc/8bhTh9rhp9OhVG9Kg4Sv+b
c7RddgdiotLacfP1yq2suHTEjcP55j1BQO5snsYLxPy7EeEP/921wNi0kt+yZvozKPR3JwOUeawA
yhAe8U/krBVkRyjF6UGPp0ZsOhNz42rItCTz0RfRfCfsBm3gUBnJ7e27Ziq7rlpx2k7+fwwmHlmR
pzOUtYxfxStUCUGPpmIbdoJXKCFyBJ8NX7NvysoN8IT1VyaZ3NWhiWh//7QSRtc21J3jLQFPpPOl
dbH5Pw8/aGGH4hDsQj8I97e458GlclA0fckLCifYahlgN5kqrxZiiB/3/vdfVL8vpRWsfVPTvGUr
V6MRLXoFlZstKU0zxqfUstIagNo8OL9MkKStBrV8q1r+i5eRZdr6+hMOayOxPm1dkH8HsXNSxANF
CfRPDMjvn91IS8JhoDQTh2rz7VdOZLm2Crgd6oo+HvEqm2dUxy3HWb1CXPEMXbEzj47N3AT6HrVy
ZJnw7gpo/IOio+6yq8LRr9sbd28fR8BqZ41FvoLqIRAsSSlDDBJ2ItI1ioNeS+2WUK0jIqxcUNIw
L3YqtnR9V9KekNUlvE2NqhO0VLh9jXKsq4H/XXU7gdFR3ExwQ978n59+nu1+fe+frT1/bGNuXLNj
NEvqDBLUCtmNrvuRNspQ0cheXNPhCWlWXNIxsjDdPPY8RlS3BrhqcCvFwb/dn4/43IEghmF3ckwh
jtLr6Kz6e3Isv4ibrUsHiMHYIAoJUbcW7Ro5+xRH3RhLSYc8qU2P7S21yO+cZzwdh/sKtyXbI9tA
sGiq2xcdDGpPSU/8nYOcVyq0l7EvOQg57xc2bGn3NKbS0P2Ob9mCOhNLdEaMrQgarTbTHqd6dsf/
AN3osHWbjm6cDRnLjvcxP4pdxCx3stSM/q7G/fWNYZNQ4YAqqc6SWt6RghZqJn/yw6xoMyuePOCM
uW0x9A1HABVEIiegjDqPP22ZfL7G5/jd0sG7Tu4gfO9pQEPHdOqqZ51inQT/ANXtDcmmkP5I+MOs
CbsqOSTHUWuoS8cHoiwpKx2LYDJco9vHfUphSw/a/YeTgaTZIIxrW/AoPyJaP8gIn3xp1SKuGdCD
7qhAQ7CXDEDATlfooSxfyca9d9DfC+UKieQ5cGIZwyUzjbgw5lEG5mQkuFU341ipxIfO05JkVAhT
rK0IWqsdLUypF4/7ynk4b7PIyDLqLXcP28OVMhHBuNacQgaoKu3+UBRRu6IdSJ6d0As2X8HdorPV
MlAcxL0lJsJuZx7Y3xbH0u9qfGrcbHJM5dh5ZyKBkqJCTazUXfnaMKN/4QsGXTXp4BxzEq7p7CnC
WyGYo4aTu7wamkEBMbQzIhVtOmAcwIzBDF68MphIg9i7ozzPPqDn0w/KKWh8uk5xbNUGUapFT4jg
S42kN7q2E1IKiYzvopYXCRZe7BCCoOaeqwh4nBMR4yQXSEZX7WGqexynucElPm1LLFLD/IWQ/c4k
tpWeJIvzDE7Bpl8P18Spy54BNlpfPCan9SnbfTftlz/2sx5uLtlOSEMjnwp+GjqYB1VLow1RxMLe
RShrDYm/euNyK5Qcg7Qgt66WLzGIqLTT4D7d3Ij0kS95W/IEF2KAk6Ol11HAR7DmTQDnOiuHNrfH
DZQlssoyGqi5CerdkvNJGIo2Ij9LNgvUvf+s4aqVSwdEQJov2uQBxZajqQove1JL+slv7uv3NodW
h2IRBFQZi3Okbl9eax+nQyb4U77BPBVnElR3QFrC4kB6tgXW+NwijuOY7MT5od6+ynY8YY+PicIs
+8xRsTGgeQf40bChc4HyGBwi5jW38UuP/yxbu97TZuwBZ71HM+fa9Pv0Y+RcTsCXiFomRFh5Lh0F
Tz9nSvfyoUqp1tzDXdOl1P25YXzkiKmLADYEJkFE9z85XkBqVtIBC1C7WD6eCM45pjHVkCnO7gck
fFBKzyOyFvJBhNxensJYu6FcY2EpSYCYeYePIrfhlMigmFjVdDwdhWbjPgxPOTT7mNPcDTV3AsVT
qkPbsWLnLxdGkWxXBzIMba1wQvzvo9CDfiBbmHiJqK6fh0jNu0UROnZ8E4sASSfunIBopGdFq+xS
cHfeQ6j3rHhHVa1sWylPDr7QVk5XxDT4EmVGvKYrv/0ByX4YDT0eg6vLmY7JJl0KCjEEvLj519iz
Xe7GMb4qcTzgPDGNjNUD8E4nHL7Z1+vW2USBtr4YRYDVkzoseUQKpPvrp9fcbqLONf1bGbprM4UY
o7NQJxD0GkcY+YNjJew+QH2DVvOsp5hq+ZnzfCHkRSSTlXj+WT7u+n9B8Y2WPuZQ4OEOClfBcCq9
mwYxYoJlgzieKo/lqL8urhlGVO8DKKW9P/QanvLGMOBj0E2lsOeB0Y/GysOjQAObaPuPmipgpGn4
y8fwLfXjeOxfV1+RRiQc3ohK4LUbvpJIo4NMppvo1eFuwR+D3R+e28VyexKGCBSdsjVT+vM7EfMi
TvBffmVkHbUhrh9QXz3s9IjJ+g1vT7gEKsWbIkZ0UUbD4AwNl6hEFTI6O/WKc99VWBVYF219qzgq
vm93BLMRronvHKLEzqjX1SGVw9ZNXzEdqjAEd+4eGV3Av26vvxpzpbQ66NmAkob6wfERANU/C84k
kgi2FACEmAAO5tRMOeq03OrvH+gssQxBfVABxQIwxNBDklHEJQ/rMqx7hboLBX/b+3JzvJRu4tdv
90QYXlmaPYTN3IF1vxPuc2QI3ImJYdTemgpjT9nbJnjmza3pCbPm2RR4pN+T/2dPJ6SGV1MioQRp
3CSWMMMYDq+r3NszjY6RVY5htidGHK5kYWGMNu5up73UK+ZJzs4z0dw3+urEVqfI5mbewXmPIh+n
dhY2onQL0PyvOt5+CI7iLvd/mS+lLiXEwmwa5ETD0CKwHER1G+f/0FcYb7oQE4DbxzyExmVG/opW
ZXD4YX21G+MErt+UU2vfZgM3IBgOftsEM8tNOtkkwGd0an8vw7d0ofXNnBhHC0xbRbYN1aB504Mq
sbM7Cl3514OtUv2lM/1htIt6v2qU/vXYmv4UCdo6R1HlgnHh0oRUoCbq81StImOsmIMdRj63S5Hu
XkMZxFxZFCs2Iw0VkUPBujgkQsYhJCONCUeWaBb4RLzpsvI9oNT5sJX2rfkycF/ipuUuL26jUekY
Ghr1d0/pel5D0t4mZx5oWDZOVIw+fS+CAUVmNT55hUmWdpKnmQlXWi9lvkcbK+Q1hIbXBd6e2H6A
t1bFV0mpsmtkkXPdudoqvvdGDp0C6U1Xeu8JExC4yczWa7y8hWMPOeHKzGOPDVWwXdi0nE4nr4eD
7VEzNJOCsPzxmgxiUSGrUwbFRHnoa8pXmcOs+xbnTGhEmFwpxSwvZTa+dQqYPI7Q1psUlgWPqjH+
lFUxXg3j7nrYWiedkFDYKjD+tUH2+T5l2S/DrIsT1bgmY94Lj10O+oONzi7xnDDAAQ301Wri5/W5
b7Yk3+AkumSc8Nz97xzlQUBWRRGF7UnXY2lc2tBSTM4Z0LkwN7Jg3WbSEL475+ohh76YUhBoy1/O
NgSUI7qxqno00h1HIKjZaHrM11frONXlMs2l2la7etl3tWVJSOkGefur7KMldZIszUjEMPE2S4ii
WNAlrTIVKVSF062S4kmzttsJRn6Y26dt6Fg8BoWIshZ2ZELmZsewOhusqVSCmVMJoAHukyQ1qQNx
Bb+AM5JyA7yATxCE/EZ3xMbDjinZzuEi1BPl+D9FFM5/aMnvKn49XuSelgw2sUnJfGqvi005+fuP
9NHeuesMQbccyEZh3KEoOK8KEUT2rIBH4jTMXG7wmooVEjCtGZ7crD5Gk+21auLJpVs+z2nugFuV
xUC5K31pigwwA4FcFISJlShFCZ+v7wfjHHHkkh1p1sfjIAHw/d/8R4F9Ie4vhSHw+okelFm9QZhU
To/eni4+m5hH+S+6cELhXNV2bnYqIaADz4Hy62DZVweTk7GEo5gpCHp/q8FPlWhysSp5/ggNRt7k
2BUGuUSY9Rxd93q/dC3t67b8ZP1evo8LPRSMpc67rzAC/tUpFitC2mdnLpn+mxVvuPwtevf07pmw
8zT/DzAQQ83py0rqSF6pM0bHsmhsUgJMUVCsmFDhulJk9RBqWae69amf0UfFRuIxvSwHo7x9lUb6
fI3BMu0LjCKMENIl47KWwIiXp56ZdAHir/NYFtAQILKw705QUTtCh3UcXNRI7yq8h6Uqa1KY1oGb
JidXrx3vOOY+w0nrcjO4vd1kTV/W57Hd+qtEpwlsvUsFK38DlaBrqJn6qvorpc2ai4SkQU6pVm8p
e80YHw4W+UKEorSSrwEQJDyYF5mzcdC3j8OnFmex4VClmESeE/FIVF+8bBtiSajXAmYZujfmZnDa
HHenSuKpAM3hDLFG6j1dGEqzGbjhJaJh3ct65cg2m35Y2aFkWhKnU+5jT1PeE/LWTUIGBLOSLX97
Uqe+8wbs/vuGYkkJTf9UuDYWtdFY3DTqX1Lak1B3bqgpUrBN86qRWK5rELPTu/oaNfKPnvRjaPkr
uC95ho0HxC+ZM/nHlamrBsNNLDdSidv5UYMboxUrxTN1Xj85l/LK6PM/U1bXnux4vxH5nzetBPi/
XnWgFvY2Y2edIo70UaBa9UfU2ujUmywnmfWHgAQCx/+xCn40tfh7vTb19I0wywnr2HQZPZamgR0a
AwzmjCvS3rtPCqb8+59bCDjBDXsUrfdJfbNDjK0IztsttzVblZxSMqE4M7iaBRy1rV25hvW4fouw
W8ui1FQAJccTYXuc50M8GdYdCijPO/1V0bWbknK/cBpGG+CyhYadvAqfKxnoA01Rb1llq8aXAAks
to+yF1U85NR41ySOW1m9LlmQZP6Qo+t2nJmt5QpK1SkuSnsyu1XCI8XhBx9EilPpiUkKiHc1cqC6
yRDwNL/2TL5Vy/9TOARRYq+vYKELiunx3O6wG+JoQETXqj4X7vcZb1rZTqEfgd1ACRYAMKGfjxLP
nhg8WPjubTEimydpijStl6+WT05jcBHXvClsZ9kMrFt3oHR8KNjiPortQa84shsq4ylENVrdWa0X
Qi+on9eqMl4MUW71cVhl4pZ2vYrzZXXgWEt4nS5IqhjhIRbcEPNrOfk17h6TUWrZtbVoYuSDbKdS
I1ewaVGAD3J3wbKky0Bmohz0XvTLtuO1KTVFJKnhwrgFACZ1Hd0rfHT5Rv9a0aJL4Zg3QsjX2MsU
7TdPhIbwjyq+uM6+U75bhMP4HLnZvRWaT1Li8KBPnI95c0O9XxHclG7kh+jgDG8x3IMLf9hMmz3j
10FU6mlgLy9awj7umYEKEtheosumDC0w0nVh4o6cmQD3530zm5ijrzS/dZNTVj6zABDCsJg5lDWC
R754HvZtj/H3DetAFS0NJel5JMGy3SpGUshJAxDMaAGp+GLcO5DkYu+VViH8ZE/WNtgPV1FUGxkg
/RdDXm9B6czFdPK9uQyhI8jd1gxrXQwITx6ssXlYp4vpL9fltEe7zo4Ki5UbNYGMlAunmBqyH+OE
g3AA48UsvIS5p0/dnUNf59/VusMhEcwPSD9LFathD5Elg53QDo+BfqACmr3U20RM8GtVIztEL3kG
lnN668RCBoahNSZt7Szb7mQUQ0GdYnq/+QDpWivx3lEZPAJrhHD4+6NKbcqdqtWPPBsFptG/XJnc
3XD9aNaNrGK5cVkl/d67DVGyI3Rp8Yq75Z0XhWSCy0SyXZnvxeoJxahKxa8fiAdqkdHMqUUCLpaX
dv1y3uw/hUymQ0II/fshZCWpFdvGvnBO4SZCyppPSfsk3gDQqY/529rFqrsPC1rA78oS1mcV7DIu
tTNKIysAnusQGjaL2Kw8cAo4NnACiM5nzDy4snqpZVkpbAVGFZi2jlCd8GD8Q3zwfMZUAG/foWRh
NOtdQzxiiFGeum0hjoHJoeyVKPMAdAOzjn7Z9W+Y7FntPItvshaE0aad13wy7lCnfI+BiQEZlxxE
GNrEhX9zt/Y88c22f1jrGemzF4GaI3w4WxtUQou9jTGdliZuUlZpVOfp9fejPfmxtgL+yolN2W9k
rKevHJHEd6YBd8NIW0P2zQFrUFSA5nCCVaWdw3EFfLko+LFseXm5IoZHBfp91Q9kAE2DWq87DPAG
6OPIuj0PGsZQqZa19KeLexll/6T7p59gc6XENfdGPvhoW3dfz/FTWrOIyMHQV0EexD3ENa/mdwCG
qHSXSJ0fbrAjdTFjWwdDgpqSaV7SruYHS/2wk7DkHhcuVSK8wZ6gDDcCM92Dmg5OUc14nryask81
m8FVNdC+5i+34WaGKxpl0WYpnM9rB7I+N3N2inttOOf6qziJIaKO8h7oXsBw4FtU4WJqyssQm0M0
84VBasKro3JjkqLhpcMAjp/+Iep66DbvBvbeXCYTTHrNcI1h70IK2gYDkF6ty4g0LjdW0HUk2mPK
LI89itmqaoxCcLNXe5Ufi8B8bnT+Sad1VTVyhP0efdomqj5U5SLS8CJmivVuFN1oJFcpexDfnoIK
uc71jgttgDynCJZ/oP2V+zFLrOyW+bLB9e8PzJ0lYrisBroBpson7QXME5H3wehTgAXTiDYeVMg/
ivonhJkO9buVUIQi9TIE5ofDNbc053BfkiPrMUL1KLDz90ZVGtkOVkgtT1HLZ1PjIOZrKvk6SCD0
27+gfDYpg/PyHicTfK2uZgurDj20JNaiGL4lgpkZvDYxebbqnGXowvCi/XhnXDNnOtY9aHqASeI+
oJIuW+8Vo8WObBALfzDhiqC64luMbQQ8yxRItzn+3hkbHrgtCcOm0pzdXzy+AAERu6g5e7IeP4dq
JpM3BXn34TeD9HoamENttJ8GDRHor2Wbzva4ExEQ9Ody2ip1JOlWmeW49XBUa1G9urWd/V/yAlb1
4Vie7DCuXmHm92WrkDtP0mr7HL3K8UdG3bClmpyL4RdAgfsiPl2Izi6egVz2okwHN3QlcDRp35ro
kMuojhE5ooM8K7MJJa/EJGoWTme4YUl0ErBTgP5L5ximAVQn5PSuYo23J+4bYCcIQMZ2poOu3H0+
6yjEz5A3BGZJYny2W0+h5Zkg3RYiaeER9O0ckk2T5EzKktn61U8VPRZWkxRMVO6aEl/Zd5W9z9l7
oVc0YutqRXAMMFgxkAF+ESf4XKiu/sJVxJaWB0t2Vc9ONWa1MeqvGNuk5G+2g5ABWFgM71JXkDnV
CZtCL9ZCVGsIbbAR4MuNaiMIRKmfZmU9rYho3heFvI1jgNHbDEYjSpOaviENroZ36NBxjUUiDAqX
cf37Xrse9a/oku8S9njxQP3mFrwUxPgF+2RS5WQG0vcm/Co6YfLpLM9wnlav7u/GAn22Dk8HvQNB
SyyodTIQjkTB2jR6zK71zy8lTrGGdQTDY9323BzvQihmhjx2GGb+dNhNuztnXx/T84j4gpPiL3Lk
9BnYumGi6vHgcAMxRtCZWd6UmER1JYW3qTVFK1h7arcaiETluDp765YF/UEgWVqsr5YyI5JdPw2m
x0s7hNL7fR2w8LywsKLmXdcFFoGeWfgPztV6ZWGhHDdKe3ih826qj+wCmFp9zo6GN36/mK8weNsR
yUGlOPr//a3T510zLzFYCdHuJmQtJHZ0iKH80uARo1N9kGvJ4Hal4SKsyNABax6leMDg6kSPqVCi
0iwtj6CLmKyAXozM7aZwOVzXdBRn05JU4LVVuXOCwu5W478doTPV6iYHgvYVJcV3oV+XH7ZhpiW1
n2mZkLP6+4CG9WEOyhXQRnAbyKn5mFlv1M6YGai8BGIvWGEi43fxf+/4s97pRZG/aSq8cWLevbe8
OvWemlCdeJ3XCfNU+WyRdRYxqtisTz3vrzf4K+/KkaWnTypKZ7BjQj2vYRtnaOvCyZFVApYRGS6H
WbLCQEBmqWwcy9VEUbexKRMmhvqK11+/6IxgjKQbVmcEKzFNPWcwftlrLnir1VLjhO6ZOXrolUeo
n16/s1pvYzUkK+fHuA9LiU0MuR1ST23r2hJR3bOkNsH/Q08f/+OPgJgKvOhrqFIFUreWzPQpiM2f
rufk7rCkHotn58ecMfTXr6D96AuzAFHov3/KZ5lc5c0Z4aynpT2H/tmop98ngCt3x1cufyp6Flaj
v6xs/0N//CpYqBvDApWMuxvjOgXmv2BHYvXB+w2cjGkzJGfo+Psju0M6TC2kzwP1ZNpYNqV7aZaj
YO1bTjsqNHjC3iGoItpeEICyjEhztYh6yklM03Xm/jccaFLpLBvg3kWepneImsxVhy+2FBWa87zj
ZVzL3BdsDaASqtYm2LpbYHxu8BucFJpAMmTYPlU/KNuIaR1bi188Sp2orsjevLSAxi7MoewABd9+
WUuqp7Kf8fdR6CMaCDS4YQf8yF9IGpdj7plPllcDHVXZP0zLsKoc+EAO04/iJ71+glErCuBxKt+s
ueQTTEEUnMnFJROrfhwBXbjlj27+dJ7ohkItwRWc7LwTlvzBn13yN4hz5x81YDrbWSgDKT+M2J8S
3VIt/Dq7rC5u1DNItK1GnxKWba+fRn35rXYGTuuW9KTJCSse1C6B7fSHgMOz3HIlz6MDU3BELUm6
6yo96O1kkbtyxhsxUA/09Q1K5+2wPuhDc4Wfg793td+GpxXFabD2S4OB8CRVzvee44ra5pMyMyWI
Kq1wbSNsjVFPncvnQQvX13+fuSdIfun/kEqQ7u1qYY7Q4n8xG1cqfNuYjJXYrnB3JVVelJUwaZNA
h/uR4xlUTwsuiOKAkXO23m6mtMdzBMz0alpWjle5omSvUPsa7oX/5aE0mOmMeRFdsMxMn3irSFJ2
rtQlaKj36X6Y/aa5SLv+ranEXrKRXFei+G5Hn5YDK4/9pyrVH8serVzw0oKItOmyqDUTs737pMU3
FGeDnGv5FQ5M36GNVaUk/VWsxgq8Z6HmY1Tc05k47FgwgE3lzCNakslpFOecLpa5+ioJYLQDrVpi
uABi+94iNVMO1FqH5xm3gd6JibRV6M+BUnuvF2fi/gjy3JzqG0uMmUGEnzgGkbOX9x2pmKF94zKZ
QfcZIvDDKryCkhki9tzsXYpCWwtWNGXN4B2dcsbMXC+h+k7Lbf/flVCvShNUK0AV9+0Fv1KmgEBs
mDJgIYPCVsg6dwY3quE2LTjLD65Sgps7yal9SClAisUcEdZDONWQG9Pg+Case+qUGeVB/FPXEkzB
QFr4FmmWMDDH4Pnwb5ckEgh+HG+LI6ktD+WoP8HoHJdkfmUcVbSdjfN/ndFSKgJbsgZHR7UIutQK
YroHUdb9bp7gV3jwCsQm09IB/HZB195QgP+ctJh4iB5dmEwcvm2S0xTlNzmKuJzY15FcVsagkVWH
1zCTNBtV8K2riobGMaa34uY7/nQnO1U0y5Sv/gnC1RDU/c94vmZ5QIdflWyVNhpPpUvYsxPWKC2Q
p72uoaLUxL6f3MkNAqSQucSC2wIydfIA0DibdrZSjGcCcSFEZ9AXNYGfRboTDrKIZzFXgvzwOxxd
3e/prM3/IfGtp9/ggfh+Fz2B90rTZaMf8NokTwb+L6+2KCGiGEH8RL1vT70DdNrep9AIeYHA8Vno
G0XbHoj/FDNMNkymeByKofzEGbDIAPex+/qx5fuo+LxFLT9UAb2CAKl0BLYLDg2RuW9GeHRt49o3
c/HJLUI5rT20Vqr7B5xNQsyI4iltxDGHMl/ytNzcQ1y9K2w8isa9Eh71TmvOCqJ1Dm017iFluz2x
Rp+zz1oRfJBV+pGykarm/1zzgcvebsM9FyCe7fHAJeI+9Pyl2x565I/Ee5kPHxaf2eDK2z8kmBYQ
7Rj9gXQzkWPPxvjr91HVodNR3r8GFd6pU2Y9eqjtVX5T5fLNRka6QJmPyyrYprirurfiz0gsm3DQ
yeDDSAAWqI3mKj7Q1zZ7RuIxsZ6sE93PBurSP7xxhz7lwOE6J6eZNnPiM0gbhpXseWwSK723DR7d
Gj547mpXn/pxysxfYgQVwCrVWTQEQrggcPDj9cMED8kh/bYOvpvBXiylqqBORGz35J8irWapVxXH
O/IYRhThY9sMF94LqF6W7ONyPDMNx9F5JdhLsXwFQ5fcAKYhEj29N+bOqYtVsZdjdz3tfcJF54Fb
cZJsfA+76062huaxaMg09yuzM4nSlGiwQplHGakLGYFtj32x218ph2YHvtedZujIrdbYwf2PYBSi
gttgpNU+aTkL8by2JiS4i3zH56xu5DHAkWYs8zDR2y8DVLlm5MXWcaGmfGYlmeAsKmy7QJJBnXPh
D2MTs7cS2Lt3pFeu5WtYg3m78919un1ajaugY6kEzn71WA8q/UWBxbUwIXd9XFuo1KD+C0QmGjqX
HxhgqXdqmUO8+rJi//rEIyKUcTxgXu8SSip8Tc26dLkJNdqOzQw0rQ7C1Uy/IOL4o2ZhmizzOtK2
KEgTkG5sAWHXDYh+wo8gkueKEWOlSA5L/yJoex+RAuvNp+JzpA3NrWurpPXQXGBWql9p6GaVsFeM
JOiaEQCGaKIv+JN1oBP3BbXDbDrmYHSm8oX++wvAG5fNm008VWpPgfMGxBIcet3hqB4QGMzo57vG
VZjpoiOtl2gAOG+VaJ5PdpKiUGRa/ch40NROevO4cl8+8YX1drjruqnIoWupEIRGWPQcmVRRF35Z
+y+MMjcRYYzas7vWN3EINLXk0iGr5Wp1RWb4R0L2ppjadpQzIIxD3TMLu90CVr00eS/tDldTbbo8
+7wHSEiUPFbnQ9foqyiYXVtff4vMvavAUfWuPM0cIjw5QRHAX+2WifYAW2KQy6ivVB/jkFpZ0iMn
Mu/CtafYT23QA7f8aajKtRKNSboRxhO4BevMjc0RmwwPm3NvGdVpFTWcNXwPx/wfp8+0zntK8vK3
jjOpSXxNPhqLeZxqKMQfZxH1SMSlWAx9Ds4Qi2tfNAfhU6y+ymOQ5LEslyX7xawU+T3uzbJWuMDY
RgIZWXelZz2DAeGTmbHT5Z9U6hB0H2U+5Shyrwlgsyt/MtbNBIXcnpUa3wcDAMSYYeJWX+MavIVN
7fpUPtBvrxV8Ee16dkn/CC6gbrz5xYWTviePDfwr5pSGuZdzEnpRd05CBlkOCnQJqC+v674gdyM2
asmdY6Lxlwv1kpzbGyC8EUL9PBCLTq5nRC+d6T6vt1mO8jYAAS+o5Q9KWq1IEAxQEeY3spyYMHEH
9N+dLH8kfwdKsMJ1IiuEIBFzm6gBMNJmCnkucCsYuPVkOTuUdk9nF0itt7SxnQxV/HXvJj1O11vD
xO0E7/uvhV5wtrCGcFEd890trEH40P7ok5LQnKwuTr4aprraVhrwy1ZeYwEqJIp5qOYW5gvqwi1D
2VgNpFMVQM6U98eV6q9xJE51F6jzRgQ1C6F9rZQPIJh+4r59xflpO+2QFHfuXBvYrlSIsbqa+/HS
cuDP0vNM6F5XlEdJJijkf1tIsiMji+z0IuIt49KbKGFu+lD5WX3zmQi6m+zp1Dib3oy3+0XePj+S
MRM2ejQIa0jMdwPj/i63P41QBbTRt8R72LxvvNFsm+uKj/Fe94EC3bbnAOVqCZcqE/eqA/eDlqhp
iyf702ONSZ+ykVaNIl6emYgXxBxPcrSc76BO0IJfO9C7c3s2HHdEgfb1xhRzljqBJrEK+66KtbM3
Tyw3W7g/inJiluya6vDMN2DOzyYWN5/UbXPvmtaZj7zs5ZuDJDFIzghVDjmUzNZuUdzIkteS9v76
8km9VgSGG3N3O6xxxRAdJUaqudjJ5F4NDEn2qr2bCVRGKwqwL1WnxREYjjbOYv0Ldi5KyjVih8Jm
odfUkl+hNpwj/SU7RIs7KvBf/f6Yx9WIopkTU6w6XlSyO33MVBwfHfcuz75tr4DglyyDrLg1du7U
uwI2EP6TyzweCx6m18XwkP4G2r/9RqkCXWZ9CcwjqYLgpxlOF0oPhKHHFE+r8qIgYq+GXRjFr149
B1bjpAqEyM501++b0krNjYf8H6H4wWCNi8H1CaX/Vi6zeQLwQfQX69YGVCTmiYIsJTKaajro6Hu5
EKKKQYecFpeMYJ2s9zHErZJbVsvAENm66zC6lRL6m/ZGyPxIDZHq6XD6gjiGG392dFnX29bUHfi3
UXPanC5zzkOpJgD22LfF9uMb1lzmNXZmGMnjma3Z9YhEdKrT7qzy0nCSrFd+0foWOtY7v0hZ20rI
aslOf082I3qF5/yVbMhV452h+dc3orjCBSskK73U72Qhm46RH1yK/mk4aE6Gy9AzSxDd5Jn8cu9m
E55jS8SewuK1QYjX141Jy2vXhWZQloM/KSb213ESXvP7QO7YASZcZr5n/weXuhDM30XYtsY3DoTO
balcibdygKXs7bXxgQgUOgKE0fxYOA9WruO1rdaeEXP1OGFCCKLUU+MpfyudxqdWNkafEkFJmhjR
LTncEfyaLY8Iee31EaDf7+OsR5kCxFLp38vVsDUoaHRqnXOPyHLkk3D5LVHTYv3GmxyCtuTZGW0q
SLANsabRrTv7WRcg0MLODZvtpSGkagPyq8R5rbPpVDfOv9VTaFEjF+gub8E81MhO/G11MfY5Lhaz
MoDPD5zi94TQIOntwMdVR1N4fZqQfMCnkDBvxYKr+BvhGvb/z28sD2vKEdxWApdiBQF+vA6awhzj
/aH2pVgUdqTE0Uz0ycG+D+3nooUOBOjpalBnsS9HTQ17H0HiJ98qFPPDzsgwadpkRaQDhN5voASh
oeAFMLAB5B0B1e0uff+mzGY8eN9KEloWfQP1K3Csq9vnduWI/glEUfGF45lFSvNR7nQBdaKrH1q9
Cn8ufwxFZigMW8PRnHpiWca8zhUeLS03QvqwPPmUkYovCwvE0Ek3XYQahkSnqyCKSPF8awNlSCpR
Ra7A88frnTeVKG7u38QvUr6sfQ4F+gzZN9DDd5QPmIO9ovq1KXk6oqDuKR0mrwrFkbCZmCjTxN2P
qTGXBeIRBrmveeWDKdb5JGoFHLMWqdtw8DNz1FCidrfh5yd/2Vm/FXg2taf+tVMxmWRlL2EyZV0S
K0FVhEPlcHh3BHDk/gQcl/RzAhFi25VXoN+pU0AOFJF3j7W47rJUPgaG5P56QH6SmE8MP6rOIJC/
F9Z+BEOdiJ7MnH+rcF7PyDLXk0auRlJ6h956wz60rIDk4zaOXv5qICqo5OXGRs4nBy0s/j+M+TCp
vGAFKtLnnadtLmnDdHqbe1gVjftrfA0cayWDK3867DrLSNAshI0nymBmUOfJb5b8GJPkOr0YyAaw
usfZyRAexc3ShITTIVwX/2o7rxN3zDePegvQvRDXSQ899May2n0neJrsXlD7EvCP7Efnk8mKag+F
RnMHhitRWNq7w1v/kPWN2bD9/69QA/sUg/owyOeKKF8ewGAQMwsTZzMbOaoIIkMmh9XyzRLLJNP3
Rx4ZhBzL3v4z9fa7DW+iyXX93yK1iDSpnw87XWygxRLQ+TFCWqVWPSe77owgYqB6pQfZKcOn6YOX
kL3a0XnLcWfXuFzG8fs+SvudrdS/8Dk74H78yeMWNhMD+RDZRjYvw8dIRC/6LKThYVmdD3U9g1/2
ugG4pmJqsfcbHFYREuITspk3s1DF71WDW4DxcjUCI63UebqRjv1Iq2FFb/sFZxhVZyUy2t9EH7fv
kUrVDqLwShVaQxa68YsWNL0QJq0et+B8yruQGBqmIDwbkfm9z71s6n83BAtFp8LIWxxINb5fol0d
gl0lF4fLSyUXcAPDLrGQNjxggfY1tKwVX2W4fRULL0YQDpUdez7a4wvHLkvSemmZLfpNXGh9pLvO
72vpPLSo1sI2L/2LqZzgq6lCPVEMsHbDLHn6b6sw6IruZLpdqJZi1N9q6WaiHBL5N1fZnPugcoIB
Mn6CoqZI1J0mDzWknNVmgGwo3BDNtqGLtgQpX1zzdCkp5agb1tRv9JLDvbxU7Fs6mIaeoZH93wZI
SpCYOTXSbdtSrRHQA7tBu2TA1eAUeJP3Pai+H3mVYhjZC6Rsc8pdOJVxJ1Xn8/coOYIi6oX4H7O3
IuCaJXpPwMWzvqk6F03zcT/0BKKsLtUmb9WPWW3pQMgIymKravpNPIcxR7Y99vYZP5C/sv5eCIXt
hgoadBRHpfYxj84t9x56/zAvLmnEpezRpHY806bBIcC9WZ149enwrPpu7HTSPW9vKZkOPQl3DbAT
Jv03E6CpHmzLW3EmLwnH3bLmva1NZ6pVdwL8E4iVQVDTZcjwTJf6xczfXCadkOndEt5mzUFGMFTc
+ZbPTiZlvfX8pykg+/uoLXU4MxZEIHPlAFQZw720wuAKLUZuOoKKk6ai/6cSeLHj58oB8JFFIC94
uDDxB5SOUdmMFLEYsBoHHZQ4wytgDUOjW3/mKurVHhylFqLY7mtK0FH7yPslOZizJMm9fOtxiC6i
/jU/HzFh2CfON/LVJTQ4jnp5+vAdvzhPEcUXMFHpSHupqgUibkIrh2B37D07zZS7d7yp5ivWMlk7
2fEU9AhjP4g4eYWDm0Zazyq1ab9LZD68W8PX3ZJIN3uobTx5sWjlzZa+/AnDPSH2qDy6/vbn62+F
YsrsozV1oAg9ITEKaSiC3ZCxloabGAo8RPSr0DlTjfdM0CUkCpC67uz6uSMFHtY8kAMTxJhwd8eT
cs7KVBXjhemBlKIhM7xIISD0c50ohucJ/cDR8vpaTv/Zsbrr+wRF9QMxXDykECLFYO27FudlnSjj
Z2Mq3+Ny/ng2WwuaKk150gLuX0z6KnRyR0lEycvsPBKW0msnxJm/q4q9nhXUmO5EQlebEE/VUgwH
Sf/xNGJCZcFd6OkaNfpeSGyvB//JKwmqD9P27fUJl8OMCy6hQ8wggvNxfgG7Lfxg9OqClToFAMqW
JinmK7Ckp/X+A6LchT3HiWd5ShIxmxoFwWKgac+YQd8d0CXVKc7rs6MKPA+6O9b8e3tC1joY/SY9
RHkOOANzTm4QtpOTFWxr8p7ha2vbRIFFxb5F1lSnn25kJx7Rd1osuoHhFkLH2r8gAoqzmUfOp7oi
spgN66CjPBXNu8M5AJx07XcyfEaL6XuwNdTmKTvb9dFQuVZsVFGDWXuOWiSZX+Q5xRQ/LiethpOo
Q/n+LhCcAnq4QDs+StLAlyzPizD3WU5zoAJWVXpD8ZMTAxqGkGt0+QXVHZWT1N0/4aHOqUrsvfV4
RumIsnRw41AzN0Pr7rkMbhzYtOUGi44jQbVa1tUDMlrheudGhBkj3+Ppovzarl3i1IpS69tmlKzt
RctxczWdfcSOZX6oP5fyP6DdjJA//nV0m+RWVLoc9myyFkgnCJ2V2XyKi2XYdEmprF7IbPzna7E2
up80qto5dXawHroKJ1FKc+ry4GBMLvkIoAQ2e9GfIqDxoBuNHHa7snAJoBZoAlLRCrUPM/oholQs
XLA4orWr5unhfVgNRBNZT+QadprFIPI5oiiEminPvogqpOWl8lvyn4Ra43Z667NbxzhHUjv6wzxa
GL/U9VtmSG4UL7eLj63F58sUQIyjlMMNxOJbWufgIqeYuSgjPqlsyI1XxbzPuY3IyODrcOzovkdg
0rJ3/LApyLADa8zhtFOPBhFpmWQR8bZ2oELPCol8j7SuRAj7wVnMdsoqgFgKxFw3nVoTa72rK6n/
/V6lzrOmZ3ZtgKK+gUmNiJ9vdADB9n5wc4gc7/dbNh4GYcMW2cqDI1/KBDvpknikDc3Y93XxHJo1
BwWEwBqiFEHLJ1O8RIGS7mzGHYNsVBrDcKsSqfJgK/+UyGQLzzVyWOvOW6bsBHAWCtqT2Q+XpIo+
fU0ZWfDmc7Y2VYvvuzAqJZq+eVJ6/GeGbshnOXQzx2v6FmXMjtO8fViuZAorhZPPEVlcljf5ZsnN
1rLCW/9bZGP1TA0z6UO1wB9VdKtieKsfUz/YGgrvbkZm0Ym3Er8A9YwKB9+ZFPKAzgGw9jlkIPSc
BwHZ7RibSqZBa6JiJ6f4Qs/F25ZyzyucSJxjN/X89Fy5qJIFFDWqt9NnUZDbTdpAMRREkJCwJAXp
8N5lrVeSgtZokfbj0G5CrBDd19alub/j0Xt6Sr1kpxrOkpa+pns4th3d8ZizuJlTeJUKJmNbuRIp
mKj6pxkB04JCbGAdarLNQQMjOp3/A/MSF7fs8oZg7aPYAM7b1rkVDf670yMchDladA1KiLoZDOsy
MMYvUwkT669AD+NveqlSxCfQvcRT0jnKihM1oBbIn7zjHG5a4nQSvXEommFcEHCUNcHEkUuS13lE
npWsO4GXFLr231db/YOFq3nc5CX+qFys482BSVf3AeOI33bHuuRDx4CyQwW0i1A9BonxBn0u1yqa
VIpUTUPZnq5bUQTwoXz2dW19TMLJefJia1CRnsgH3bDV2yI9dP8cpFK3JtE0f1A243a0Hzilawvv
7f1wCo40Dv89/jVHbzhpUIqxb7lirr/f65jGo/0F33sIA/dR86LYjcKlgSBHiW86W0Y4aIcVL/UT
rr939F8uvID8Axkkcv4rZcnnPCpJgvVgJToavrowe/NBE1l5n3gyrVkgj4Dp1MAV1opMH/0ZPAoe
gmGbkz2gwPct0aNB4rXGppiiFXxl/3HvVJDGxQ8wZgYAHxSzRDaWIQ6QNZqdH2OvEkWEs/uVFy/C
K0+yLmLXwm9LZ065RMC+TlNuYwo4u1UTf6fUIaNaY7bXltlTBBQOCdH7gSZhaRNxfma6HjN05ljU
Q+y6pjTVyO2OE/eQ5LrEZ9YIhBtROU4/FNdKUiYsGssudjnnqT0EHzInoWrTCZkjh1YKJ6AZ0h5/
o5QKbPrv47SAcHcSTIy+BgrjPHBEV0pWG91jKWJ3Jjz3/PpQJgo+iJKt8osbZBniES1ITofQagIj
hx52PpHoB0QcP1Wf+QD0ewMKImLFR3VWNQ/ppH+eXizKAopIfCz38uKLiZjeCSWDvp5WwyS9kd5b
xZHIaDTBDMsPdloitgc3dPHh0VhxBJ3lBO0Y0zOTrutQ15J9OnhiZA8Na7f89TQOtYUgKiULxh4U
hxMTkozvYS3n6i66me9WEivhxMm7foBSXarLD/9XrWHzqZRl/6Jq1WZGOT7B+gWATbohSjhRmplx
qLi3II7clMW2iv9f6xnEAfAsyHyBsZYwRlSLWETyBVGycFOerYo6c2PhSZ5Jtg80tX8gI9p4ZizH
RnQz8L6NpJm1RlVek84bVq85Spv3ddH+tPzUQeuIgJxSjCANgEoPfLNaniNLWdCtt59XX+2xGhq3
aXICBDiA3xKEw4j9QRaw19BtMDcLP8wQ7NNU+CDiEsK4mU3vGidaaX/jFzictL1U2dj6IJBF1dJU
N7NX2Hp8dq5Xb1ZPMfp99NJ3bTiHS+k6a7IxDJwzPSrJImVcxYFyWRfQAl+Qql65PPcL1mi3T0VX
xLrcXH/vPCopy+JjkQ/9Cx8ijeaKGaE1PYjESuNLiondBY6qmPg2UCmKH9ywc/MZMZtL+T1tI15C
jzcia2t13e7gQ0QtircNquzB3e6uMCq+vZlKqU5Bv8ElVHZDaRbLTo5MTUPzBC3QqzibO3yup2jr
SfHe+rQO4ALFVyJLLzL0/bS1pLsm0p9J+msjevfE97X4HLhOlliS+TqEWtRiaC/sMYmpxJuSpdG2
jrpn6zNZW2HGG550LYAxttNlKRMBL8/ZcCVnz1LrT1Nr0QwkNGNfzfl4YT8xDzI2/536gRozNmA0
Pyy3/qABsuPvazgt78/TxZOHPTqujWaqwhQdZJKH+8owFX3qcDQuVy92m+SI+dWmQHzBTsAK7NKd
+CoHI1z4XuaBOxNPnwdcuKgE7wH2Q0OQi9zmvFobKA7FcKIQW1/IUhUkmOQpiIsEwfHixVmLSJ8Y
acX61yeZSWfsODJAA/fGKOyV0ij+voHHNqohlnoKkLfuMglkyoXzbpimNKEZx263yrepl14JwRko
8J3hEd2PqR7ZOgkaagyVWBgmpgSqrAWY29gSuNu/76Km9HwZrQKYxzRyBW8vw2ulmqCLsBkJfqeW
QbP3MlZsFFTLhsveYEdnZSpZMmfc99ZnRkCkKKVEoy2VquNRh3b968Bih/Z2xk1s0OmMWPFDrJUa
zWC8SLwkCgReppAMVQ6oL16VPaKv+QKU/nM1P+hHSO0XrTNRrlvJW05bI5Xj8Tg28oL2kH49YHCn
fcVHryJxcQn5rHNw/0mJ52QMXrizKH8k3TicZNMgFOHcdcA2wbVTQv1gUvLr7WKZlMAuiTenU7kQ
modLRlM03yhquWIYyKyEJ10tZatFUXgG6kZvjTeDLvXRyqQMZh2WfPB4b85UlWLWqIKLZcKalBhm
Y9zH2LygwqPSE6n3hJk3xMbeBCUE2y3fvYDtYpj+13sfBcxBDD22p/mZtuUJQpepaqoXP+TLM5xZ
goXc/YHVL6fjdNcuuwGnekf+u6iq1geJDV3rwfHUFiW7yCKMzNNC1nURD9Q2IdXuFMI6zWtSJx9l
mjqEabsMSepd/vbvvtr7eLRaqJKKcqyoRxrRtZ+HQKjpn/v/bgNisKKZHbNrQDwz0OPqO8UaTpAt
gURWu9NPtkz/SrI10P6qh6iI15ATPIlBGzGc7EVhT3R52/KKGcS/oZ3vBwzwLrQubdktWjE2kNxo
zdgyO7vOfRZoNeoc8zQPX0gtWKFfEFrtbJEbDSIH+6X6rhNHj4I8iiKIoWPaolysZwK8wNOznJFV
Tx6FakFMfjImtPysyo/zc1/oF1YSLSVCc1UhwZgv/r7PMDGgDKSXrSp1FvYzJdCj8MNCC3U/uQW7
NowbGmPorO/OPkMC0ktkjsHyZ3oJZHDAMhYBlGfdg1VtmXxMoNAn655qvGxJGd1MFS63HW8iDeGz
WhtvWTAbn3x6jzgpa+kaOp75YvINj5+VzrIhc49ZTJcUPdlkmIn7BBv48DHpxGWoHUNZpSk9U98Z
+UWHONUi4OAVOdy+QV1hh22euqrb+BaI2Nvdx0fUfg3K+AOu68P3ISOWIdvzGH67At/GF9e4s3WC
h1Fmh1ZdxQUl2nr8tqOrUb4wi/7euU/PAeP5V7bCjWecKyInFw/kRrYWGKJmSWVmewFWfPxQtn22
h4o2nPqE0Y48xVdSAab6f9YF6IeH3xXY2JDP1H8QeNr4ustTcnUmtWV5t+egEZRQPODKG0+hExZ1
pjm7poMHQgmBZguw3R2cDbIMWy0VbKgOhNtMlJKNUWGrDYVzi3EBLWZUx466TAwVRC+1tOA/uDje
1+eZ9YxLtF3647+6pgwFnAXAFWgwaethWXExrPPg7hA4eDrpVCsd1UEYyP3R5cXhEegPQNh9KG8H
DjpPocDsQON33CHXGAnYpAc0+QKUMu7Qzs8OEZ22ej85UzJ45PYlh+nJaiNY6H1tmbCGfX4Klw+t
eVZI4NWPV9uoNOGXKMSJeQDGodpqvXQ3YBpFcdvdIT63UrVOd3nfYHvQVlHYNBjNSTSXelVpnqI1
gOUElTkJI5wu9RqUwmqp7YB/cXYWJmn50/Qwm22SP1t9iRyB9k2M5sQrp/viLumVKViPrP5Qt3+z
S5pRhHLyR54ySWfGbSKp2LGBpqStJAMr2ZWWTHOJlOWHBonPXgjnP3WaEBD4thOWb4mR5Ge+VFfi
Xbycqa5P83hSMGXO4zTzt1H951vMX92sTSJZdkA5RWGUVSiYx5ONr4/spQMNKPJeWSRmCy6YhWDy
fHRDSAQigfAb87S6kOAZM/H9v0gF4RAt+dDvL3gZWd5a8aBgEfmGc+7mJAMSWHpSnrc8rstXwcXn
P2a5Ok078viMync8xdQb824H6I0mVvkl+7kmDrTA1dg4891U0CBoaFUGEf56J5JG/CWXV4MTzfHu
JO8skdQwmWPaDT2aFiSHGVRG6P/ERpGj0cE9U//3wxbawb6TqInqQs+Z1/floVClEi3zgWDPzLXb
D1QobnGqRX/C8fzLWVQLNOyu7tXBA+zOUgntORwhMWhyvDmQUZQDhK4rLTcv8WoMCqNqe4ULgIXD
fBfL5XlfJhC1mbZAwYpSfEdCPaUTjYtmGaYzWBFVRHhGRcJBD0t8l/mHchKzk5vLNoSs834DOlxI
oCwyytKOynqJaS1Lfg/IBLdtazzf9ShIycSCwOzbjOOcyYlonbMkx3sVQcQReRuafXHBtl+5WX73
9Gz8ceEuGh5g2qyFI9LdOdNZMHQWKWQQltv2WtFtQ5JRyhpVsch/6h+KSwxBX3Pc03rFcsjT2xks
OUB7ZZsxCbEGYTCpQdg70FrhAcqzmtBMw3hxutwnQQ4UwketD2cL18efqmzDong/kGdeIhW1FtS0
AN0FTaPkFCXsdy67npulVpDSz8eXRLJhtHecXAWCeUJrRBSVPxEWVuFgLfrgTRt4P/P8W5yrRi3F
BXxkTx4w+JsvxDN/dNzB3Dmlude/qt+HczZUL2PBhO+lVV3FHgLrCo/0Kh3APwghHWAk+tvuXWY3
4IIZWc/kaLHS1PC3VDQaWZTyPiFgzIT7JaHGuiayKFh7884oMCUeBeMrTcJiz60+JJxz6Y0VOkZ8
odkdl27TBMoIqtt+xrGSdhzl13Cjcz5x/TwVDEdvN/pDstg0VZNiV/2q5mxAuMiRcr/aXZFDHXf7
y09FR8zLKHQydV+6AFQMyiXUpkyYH89OtUgp1Yx/ncya1Uoqrz1BK1eX4Wjb+oBRrRQ9NMwVETGk
LS/pExLCIJKm9JaIUpvd8B1Uuw1IFxljL3zJBNk6WNWJpRmELA7FL8CxU5epi6s2Z8RIRV5ZtKUV
ikdPpfcO8aHk2qhjrHXo4TtFJQpIT0cnz++Jli5sb+R1smZr/bDtFvvc7+t4Isv6sLXKjqsOSEUr
aeQqg2XJRC0+bO1iBP9NDUK2lPJNPYcd05uJt+yioPoWWvBz867LS0ER4Oxry9aumpSbFaWx09CZ
h4LPyo1strqysAEtA4Bvd34oLjxCgeU3USVSJWdIglEHtSVFDT108bzYh/c9jha0UCEc0sH/vgnd
OC+hCfkfKQSb/D4N94rILD+eF3FxSeGChU2E9w+/f7dpoG+HzjaVkmrGctGn8ex0r75Sk8cfSO4E
a9NIsYKceiyZums4gbhFp0q/oH94e+XcZY0T9Nj/NnVJK5A6zrTlzNra3QBzsaeYqIpSU/U6wcKN
8nw4nF2PfHAh/dH88TJcnPiEOkOSpagUWgBNqGA3x1cTBFfzNh/kcVRbIVUTOwIwsoosvMmymiEy
VSKzZvMfSMXD6wds+siNeqD8VmN0ucX64WkTl79SKXNmbKmRzQAVtC6CCd+iNM18T4rbPUIRPUQX
HjHVIjI5+1vMyzqvayBqtsfrXJzu0nTxejxRwySNYGJZnhvfYwysVNq6gVCvr+6Kv8ZQbZMJGxz1
k+wzEvOumC4u0ShK3EnzMt3wobf8ONSEcuILWp9SA7gCJk2DM2Ax2G/AqJ5wDMtYKfG3Oxp+Fssy
y4bDAUyVbFmaRqgUa1akemvU0CSBpoBkM0i+LJrHDbbIU8AZYOuPVZCDqJc1tiWfr/uYUPu/fie8
JxzIh8B2TJpYImO4ePZTwGuD9E9XomCcrkXqoWRV7xQ7+obzrYI91mfj80cTgDCRZtwF2c+9XhjR
9VDwH0EfdhYRdfBtOKfWPNIYcrfQLyLyPalW/dTpxoyxPGdC3+73kjyAyAQilSl9PrTggJ1HPkii
056fErwPYQhnBpJZtE1zwb9EC+BNSve/MpRRECR34kTgqtR9BOkdGpfnLZKruAv2Wl9RFl2AYPIB
xTrETLsGYdKNpiu++2tWNe2+oPoySCUhC8Am5O5uZ9l62jZMbTmEtaT8zGP5G1kWCbH2MCzz/c0i
p/m/mO3uWxVu5w+RIOpwWkAiV0geW7pjvycNwoKegV6jkhkwM6ygOEIO0Jg8us1HZzanhcH/RJpk
WTlQ3ea2oGfhwJfYWXNUApR5wp1Hzm4lrF3Y/knDPMTSHQF/oeY+8ZATnNuTaEmXAe2EUDT6ewSg
hW1t/tL2qknh33MLkRX/lvKu5wZpoot1Jr4P1uUIz92uzueGCSyFgcTPDM5ttlGfNNEQJ2P4egkQ
BkBoVh+b6PFiSOBFjf3O6gntPI16Eml8KiZLdg6Z1t8kyHmw2nOgQxCTfV1j/MZcqJca+bm1Cgyo
Aqu/Tgs9kPA8SuRNc2OptInByPl9GrVRLZlRJuKRpMx1KX8FSqobpHIceO4Xn7MdFqb18E1Two8D
4uWkcEnwc2WpBBR/AA8707W9sHHej8N3mCCxd51tAmd4KwI4VI1XKN4TfwzGYejIpDAlULZlmarm
3EGzJ8BjFVRQmte+ljFyh3DvQ2iiE3HP34eNUIJ2wYsoC6XoF+CUSSqPLEdLdr2CElojwXy+uu7a
mZjoL7+T5svJpbBPWffwrRbFLFSOBGRrZA1/iQn0CF+u/bfRuqpjRNBXYZBTY4efPTliTp7QNkIR
TRm5WQMZI8TA0nU+W55yqjqxgILq31cT1th5Rvgkm7XuLaMJzZs17HzNDVUsuiaC4Lv36JWPsPuI
uZ6dkbtdHN9qXMKXfAQe6w/cDbBgYg4gqe2Av3cJIWHM/KdchMVea99b6mWfHNJxE3mrwMD4cJSU
/h0cen/ar/kCg2qdO659THiWNf+kfkNku1HTo+5jBE/Ek8xJSafNB/XqcRh4sLh3H4dyQ6SgUsd+
NHAbzvtCyCjrdSk2bINP6BnLipNSdJzYxXYnUG31YemlmJ3gk8egAr/ZNk3m6K5Sax1mygY+K3o2
FnQXhwG1JL71DCE8tQBiv233LhwSukxMc1XVG7F/57W3197KkzVHhVOwsjfy4zg5NESN889qfBu9
xt6IqFGDS+YtDGTLuANVHKAd9N+BIM+hsX3SkpNuAQw3ZzzlG4jd+95NFFOk/oGgVTh1nbozDYX1
pCFhayE4jMrnN9cYlK/J/CZYf8X6FCo0Enm4MrdXEPLbs+5/LEtLlUbwWEIXHjeW9HONvdxrgnqX
Be0vMxujangAa+Mtk69xOYSPfKChI3r55/HsDeRd5PQxNKNZfJHG4Itl+F7/4xxzzuUCEdoq0Daj
kv/fijhi3ARxN48Xl850Y+NbGqZDf/UtqTWsi1NDPUyZjriGrAH+h1SJyd7dUwrcFjbJFv9EOw/L
criYFg6mEAcGCccErZjDZdaSnZiztekDkXdhTY5fM5Pf/m7ffZoNO5tDEItvfyWgQTp2phHYJTYW
SCPGj8elaQIA2ToeNk4mliwQrW/mwGikvl0+QECyAq5FPVvSHDTAUqwgFotHhXYniPcT7YrqhrqY
BceiKBNGBlPdysEGa4yZ5Wh8xcAcvzeQPztNxhSDiSDMyIHl+ILoZw4Mn40YqObyRrgL1UwQK+Fm
+gIa/8JIB4ZOFTdyenB++fn95g2NhdvzuKnZvt8IWKqv4qTzv8TMWRh5qNBHIG10xM7eQLbHHuYH
C6We+PshP2utbpn+3wFRYDkQtGRU3FfPFYtI70lMFr9e+/Ev+RaDO3QxcKjl6eVwZs7Obo1S15NW
mhjEXE7el9hB1/gDNEPmeMrn9qhN4ICa7Ned6xO1NE4f/Qomw3oW1ILVsGDCUwBgM2TjxiQIz98B
xNlnWgMpEKG9dEHRfciUm4spA0JHBdJfYpGu2fJYY9bwiioM9FCtofgDsaoIV1gDMQ4z+bs0FEfy
OVfgMCwzPs7QV1s+kezwGifDObbc0fruniS5DnYtc+jo9EWGAL/qZk09kNGPYqNhshpZSN6aCeNz
8bGGqQ1NQbORaibcpQvEBMN0C/98JSlaUEJkMICmvNerphcqtSP3zRJrbVp2epznfxuDvkMg4eL2
OTwsg9sg3TyshZOvyj5/mTUwCHuNbqs6za6Sf3/wPpEAtDK9WGAy+aPm2EIQEBkrlZkuPAIM1JVk
63E1BGUBnaRgYfLrjCpxjIt+VyLGf8nLqa2UpelApY25KAqO9gykqwdCnHnOm4qDiQsj3fsCNgD6
sqFqehGH9ymjhvHEZvhWD+ht07Q3hW6OYJUbetqpeaSUmnopDbpW+sJEfwtnl9EdzGSQfT47JfRH
MekpJx53AoXnoslJOa8MVk+nKAT5mf322REiFwEjzeeopyIbKiSdx4+eN+nJyms4ehgZOWEb0KZD
9a0151ujl8lgX+a6L412AMPbF0Bu9yJptHrnLnLZ1NoNELDquU1jdyZNMDNyTgVUY9a68EEgjw7I
fq2d4SWiCt5J/CsKw5u1BraR5UMOxNxc2jQxtarXnAMQHYJyLEHx0pw6j7QJK6SJ95bOlzSemIku
mkfETo2t2/IXF6CFZerke5INcM86pnbACyf+dg/RX+jTi9xqBAY5lbVjTn5czTZUPRhONc4YXCBz
rlIV07VxoJfK/dkgVhWrU6/DgkHTNIBotcbIB4HpGe09Gdf+kqBqeaxmwZkN6eZGT/8uvhU15/nH
JM7asz+N8fICZ9b49yvnMRxhpWKdV5GN6F4HvWvj89EQl84knNGvTQ0pKyTQtikKRNyDD5zWImy2
p0GferQ+4C6e+jOemN5qOmZEW8IROBaDvYC743v5BbLwZMdo9g5qnpirMaM2OCP875UH9s9hY8jc
OwAyBOMorhqgs3CoBalaWwc5iZ7Ub/uKv6Qr2P9EOrNQvliKV0YZfGDw57E237lSK/zV0dPilPUg
iXVcp5Vp67SDmzQtXeMS8eB+oNL4c4suIh7I0HBLqzh8EDKgqxl224unW4xrF+eZwB01Hnpp7MOX
pibsanp3U02wXMk0AwvrVfW8Tho48wiSJiJYilDLZ16wg2expFCuzKqtdBITFkAQBspWsQlMT/XL
LsCrGodTSiV8CHqorqJ4VTVDREOFS/UbDYoLiDh+36IJu4fUX2I6QPNz9mhnsDUyuFAkjiWKJpZk
SYNhxYm5UdgKRq8PFGhrwDXFYdwAbB1njsoDdpJYpXBysxTRY7WCXRIY+Z4+vbbYMr/OzdjfvGMz
jSZbyCHqLa9G5uPbZEejFJVqQEzpdQPkpfdIkmoJECO2tq0iu4wdm/neeTq/KJMgDMqPOG8//dVy
Nzv1jkHMFqbiSRNGq5y6S6CKQ49OrMF9eUYS/Yy4lpCjSVyeb24h7rEl2dAsrVk1P+mLFd4jr2tc
yxYvIwCqz1WFz0R0WPbtBl30fMc4FDuTWr4MsjoBkS1USsMEfcu1s4+0H+PI40dx8S7CSoCtFSqW
J4sCu/joj9CIiYR9ZYJlXXJYomKipc8KT9PRlaevuzYgegXduU5kVsOMSoZhu09qZao+bvz/X2lL
hPk3kDaCqCYGNekOb4Eey/iva//h8NDhdlKL7cd42dOnVTe0Cg8DjlIffoIWv0pKuppcKUT7MBQ0
q+d9zdzfDfxu2INoYrs+YwKI+v9PU/KLcnZ4jztBswFIcBGjXJnDVQekV1S9T6asNjVvk2/ARLdJ
ZxgSzFCyve9j1oXCSbgjyJ5Oj0XAhtcwk8k6E3iRT8EhlP/5b5tn28BxtRgNCqoXw6Qihj6p7wTn
Jsvypi/u9bikONmd+aaY6nIPDO1qHRS5yzwGh8YwNeD9B4gwXZkMy8Pn56/WmKhFVhQZiIbkt/Cx
YDr20lTDw/DrlfwXXER024knS0N/rB3S9jkCNc5g0cx81Qzc5Wsf8RNenR6Ts5YN7eWv8KEKsm2z
Ymuxf0QhuzFcif3siMVBM6/8IzhGGmMCKA3/bFjuimtKchvDzcKJK07qnNZnKXBC6OIr7ez5kx7W
pxDY6jVnDdZGkKEJNfd8lp1mhBmhDpQDEFu6A+6+0Xmydg6lpQOdVmct+4kJVGCF1E8At4pB7fx/
kNWuIV7LD5pjgkNWqHqMYBsmmOe8yq+XMFGlYVg+/bAL+cH3KzoLgCcgbJk1fqO7lH7tpKnDMfF0
v0XKhJ9ndsiXcdb1J04KT88tlhCwCabMRbcmcQT3xmK9zq83mIiUp4gYYI0CG/A/weiqq46ufyJ4
wr0K64BlqslQh+22mj6zaLZTNzz6GGDZ6l2KQXqLyBTPZQPTF/Om4/n2dDfTUXmbEec9g4Ot79BA
8VtLvNugjhwzdGliiciYSSQK+yoK5F3WhDVptahwciLncCAF0dTQubtiJzZhbRBtvAMWvyDYcNCk
81bBcVhOz2opefzNJ+YnKvsoLA8DzRoAeRcIkRLy1fU3hEmJEM9oX/4DCjl5UE49/aZiFPi/wuIc
vbLNbz0IqkAOA7XTDlVydRMMb7zrNhn2UQrfU5x1m/1pZZwVz+KtowwCH3UQZ+YKwltwIggFfYc+
67mX5F87RLXl+L/vPMhhTQd3zh3xiZAqLivxTL67Zal8IT3nSAr1ESyAMx4D05NpR7Y1vSsSRaxY
lf3psEb1IvhrzpYrFaPyoSZsIA4rywpQZQdeLigzb2lmGYXbgT6vjUPbCc7bLDIy2zvCLWolQ0d+
MCPpxPADvLMyM8EUIPoM5vMr6VKlMhe3qIqcpWVPNxaAJEo4vady6snubaEcv4RWxB1MDeoTpYF0
5y+XaZbmVN9yt2aoy1W7Uawo2lpi8bxMXk/kB3wNT+cUpmJXmMSfJf6ANz06xw1rRFgRS5CwcatK
EWtQdy5cvXhcrf4OC8u7Rw6klqxAqlFA4dMVsZfm+mS0aO9HNihwWbxZ2z05418vI0RM8A/dSnCs
h3lx9CwyBnGbyO4AZ4BV+DWTknIJHnDKlyCWPtx2AuuaPHKgXiEerz0ZTPLGDyDnCKocFzYX11dQ
pQ4H5/oATibTldaWakfJLCECpPmAT81RmcGUKI26W9i0EDWKD+IiHDNLvfylvsptBPvCEPxIqDwi
1btfvcIi3oqhmcUODnRlS6jMFPsgwwUxzxOA/Zo9Z1e6dE7Keo0oi3YRwSRB4NXM2CjUdGtkp/fi
ywhdN5aR1vRc+nnLXhPoucfBYkHkZnY+kOAECZ3iKs6kVnxYhRnp/z4xEjmFwBpezbOaDoKByR72
GZTiQG92I4w5X5EQ+Jzi6l2lRPIf0j9XZQixzO+r5mDBvmxTjCa6JVfl8mXnnIu7At5ex53QpsHq
5OokW/pis4SHP1pNVvIOPPBuxrFz9gLg5ItNsuXdVd5SSCXk4Bb87T416NnopAmHZitOHRSI6BtO
hXkGwNUpmHapl582H4/pf6TyG2Hzo6PfLhFymTOkEqc9M/nyA0/dYcH9gNwVA7DvZG+Y5Aez9pNU
FA3tEzczPoX441FfJ4hQk22zaEC4ZmbnQOxYcBrjLrB99ndO39BPi1uuhk2VseBrMGz8Dzijiyms
eCU0wstqu2n9XHLt32XDO53j8DTG3/zh34cg4QB2xIuR+znVz3RtBF3iiv9XM6iSs0QJLphc4+MD
exuPFCgjKWQkt0lWslUx002xK8AsozEE5H8xk41hoLoWHzCCfnSmvHRlSxY9oAz3RuYihBgDG+KJ
w3Q9diCz8tI61BZC+N7kx9XSpbGRR91W+KS/rL1WwPMq4UKN+CxNSC3XF5hXl66Ufs+5rVS4mEXL
DbbtT817nK7hUY8GkwPxUiZeTHrEpibvymiiEurjXAxX414ifEe3h2mX6pfYtFMt2QIKCzphJ3Oj
JDRXFyqYBntx+Qp1cOqS8yoED3QyHtsf6Neg4aM/aLv1Oqn+PGdnirYS1wJo1daPA2LeNY0B7tSY
OtvgB2vaOY+CWF0pgYCmFb5GU4sko1D+hZ89k+xBkkNRGjfykKaeE+wgz/C9HT6jgkHpQ6qbdRvf
hONzuyjT6025f1Fj6i+nTgsqLvBn1QGXdo9gE9alqF4o8wfvxq0GIdzGT9wDs8cqVmHaU/JMNJeO
D/GC7x2EcYU7c+iem2S/BTMmJBpacaYR79jX+qVL7auNH/DM+YhXkqLm8SYfzcxfsr9Wg99Jtfr/
AtNyPQHDVbwqUHSN0wj8GqgEgIsoNRd7fmWyyfbOGjNx2ToH9VocxakSVyx+fypIqB9eqIM5cRYL
zvoPrcfZ6vCuCjHzmrqt5bb0dKmyyRaqJ6P7PPFiOGAQ3qUg1HCNHb0IfIJ4csnZKk350lW5msFa
N7vUNEuMi3t7Y7Gr9VhOwI+mnmXFPrPAxaV0LcM55rri7yFgokWOqfl2cDlw/OmDw7oRpWOCeYvH
kv5zg2N/9aUPi5M+kzlyKqRd/F0jrVYAsJ9R4l/nmk8zS81AOGeslfclZzTOoLsisB0ST6iGv6rs
9fZTGqb7GD8GjK+O89mH5IsSIGjg5jI8lSAGSlCmg1+fbCZZrTKd7rxVwl7gIiuG1oA25w2g88/l
6/mipW76JX/Rc7V0xtwUu+ZipZ1txh3Q8+X9GRaAhCCQycEdbVlCLIrQSO6WkGvMaHO9VkOTAk1S
lJlLoGVSoGzRADuEAv1M8MzOTUHIPf3pZKlfM7gr40/AXsmCtl8nBDw78SW94VCuUSZjuhZsPRtJ
1maWPkU17NmnPy0iWNmBKDQaBXR1ydmqaw1OGiK3psMRplR0o57m+Y7Npd80QhihdqECv70mk2/A
G65yRavJ3mt6sywh/K+11B/6Ukr3VdYwCXyq71oJnmQRqkJbvF8/xPC0Q1tLbsnv7hxf+TXQIDV0
npfWjeSMKQKPgZINt+LSzI537DwQlfsyeKuks+tF1bCh72/EnCC92B+WdXbvODJDSwQx2SBK3PzG
1GcfgV1OOBnyL9KvVxD/xqBYQdSJ//M7qL2Efrym90WONAYZa5HWr5yUHfGE8R3EgedS/Pre4H+W
LLaufpMq4IiPLrRWwuejTHPlUmy06o0nPX7+ifHh/0sIqfWigBWqmrdos9UmQ2Zasd5+T39p+E37
vmArIRo/tKUGqg5OB/hKjH49442WyXqjjED8deVaIb5eHyjyx6Efy/9iM6VwSpRvnt/0cWwG2FDy
UY+nDIgpjZlrHYLQuUU9pQwUl6k1nkZc6b5I+Z66PFHu0Nhda0L/A/ldw65pgGcX3I/kuMxy/c1D
XAMrwnQuHaS6afp2ZcrNrKScEoN/L9LNTV2KgpT+WKiRG+x4JODmwuInQYDXSIRG1P/PBcPqsuK7
1K66vmtYm6p74LAewbz79DhnoiKM2rej+0egBWmGXDTD8AplvpPkFaJrCStAturzpspaUNQjuTb7
XdizpTcI8+GxGy6RKuTqNqYmeBTS/24opJ7LhTqA7d4PLWHHh79ejMNwhstCyPI0c1p1DpmpCkCT
LP5ekkLUBQe32TFN4QrNK5o+3rjos1x+29+yySCUnpAHOEheKcaqYzLpgi2/Q7IIeJ9fKS45ofjS
XwrHMVPZW5yP6y/i35z2qZC6datZ6VjuSWhyDCmrGov9kAuUPl2cyhd4tQCx/1+QVuPUd5+uULN6
C00rq+VPzv6ZBdAUhz1vdxkdR+dUH+ufslKRgiktLrdzOdL4ZkmrRWcVifauKXNehLFaH2m+j2jn
Cd1WxAAbOIVt1vjNsRZYxEl+aQLg0oOu4gsYSy4sOV8GUYjass2qNu8lc825Et3MZjBS15yVnjS1
2H6rps5T7QuMo+RPZaeZaU+N+f7LrX17+AwE/LXw7V3ti71OYngBqwO9+W2dmAdsTcdXEdnUfeZW
3Tf7kEch/N45tr9muk2MPFnrp8w5zaJ2ngUJdDF2RTRj6U65/tHF/dYE7x18gky39m2pxSpec2YW
B6S1DGooHUA1RBwNQIu+CO1hCfcKS8UD0NK5KqjtCAjBvFzhqi8ZclTGmGB15WROTLTMATTksmW+
fnGRDgBMEVMl76SzVpCaFRyivbjt/tSQ4q3YhxBKzE2OiLvFlSr2KfI6GWNjG/TzYTpmEkwBz1IC
2rP0OjpmnVS+0Ucw8KZsryZVYHKkd+YPeqjM6Zrrk0MDpoQMLoKc/fsnbPc8K4+KIuPyyTON3oMN
JfUAVIQBHbQaMSyTGO0AwrxmweUjEuX+BXPmE1T3oh1YR4tHCV0TrCOy34Ox2mB7r89+pHzEe6ry
uOo4MnFoczpACfQSuPWzwSfnsBwt66YL9LFTGf9TA33nls3c3YGbenyvIc0xay+oPIA3sy4AkWBS
0J5wNq22nOqK4nMkbYGp5HO+V5ktfukQe4EEdXWT45b0Fl5ZDgW1f5+rCJfqMMScHCIm64VhM9op
pGT9oFKIb+y1r/3EvuN/U9wZK//wjdThSUh6mNt5Xa401e5sQWWDbyU0B4mlHyjYTZJDtXEGuEnh
xdv3GOzj0VBN5bbFTNoHjAZ97UmJVX54lSXbjcPHy2Eu328XCWveTAG9YYfyE5mPSV6FZdhLw90I
T4/Z0Z44RE1he8uwc0XXGDCVUdTeqt/b0UVTtBoW7mVml0ZKWmAVUWCuVFOI7hA175Lj8Bjkd2Mn
SVml7hBgXChDuQQIreUv8FDSm/EnL/WhxG0RBdQzjmVlKDJ2RoQ5beM782ycbnB8cJxTS7e6GmN0
vTDTrtO7BjKtl4GfX0hfexlkIrwr0h21oamRDgaQyDGHXlWfR+twaRlmIdcFlAX/FpmSgT6EeWBJ
hYTxME0fz8ktjDuJfT+IJSw3/D3/40E0s3thLFQ0h0oTnIdyYpiUEAcO/cbGrSDtoZAjTCE2uVzf
6+H6KYhWLL59N6uTMU6r9JJuvUV6QQAM2ljNeXLR9OIReD5dTCC9X/KniQt725x24P2tuF9zC5+2
Dn3ynm0Wqe7phYIrA6Ea6v2l1p6INhZGBnPeQDZEmrKmZNufAILkYDHPQHOqHLYcG61wUEkgLypO
hPOCFLfmq5WTevXxf/GjRSZM8JZ3hCVlWDkq3fuPlS4FeGbNb7Efc+pWruINblriwtSzSGm24jo4
TV5uLmi12SWkegv1FYAssKhYw0wgFAb/ezOyX/lHi3AL+O6LkMGX2xnSFjBGAI3jhJ1hZwm+DXFV
djRUy4wo6lJdQAHy2cOknpOFUabz3/gmeik6CprEVR/xDUtQH8EhR+FlgZftzLbkF+h01UmcWImK
d8uZDTBhTBMGXJdn2Movp9qOrcphWTcF5A9+lWeF4J3AArJB9mVDO2Iep4lXm0Hax4YkPFPm/a45
o3TsEq+1zaWAZu3J8S4RuF4/y/oUSS+vHedwCXcV3lkhf8kZ70snxOkfkQTXQ++tcL+f7nPsE0b3
8k4jFwSFhuNF9BQ/4n7154gZjVqZCzPRRExTcDH+gUw2NpB8j9ys/do9WBE3JPdi6pZu3DEVUIuu
hOO/K7O58PENuiW/3Cpa88uqHVVD23kK+hbVVxpSpSSA5H9DRuI4hCM2Z/fBsj6FY4+Rg4F6/zP1
DITxm4PTjMzmoi/R4kzMu+vjggo7yIdlOA91qNUaABe5cFK6PSck4fFeTz7mghzllbsSTERfg8Zv
FSzGY6bGOsVMzMKURwuDOWL/PEiRObIT0BbOKWMwbCZXlRntMmysC+h0eJJbspMqfZmeidDWbIvx
oki67JuJIBwb92HkIFRH53T9uVvvqBAkrZ52JoHlFo9wyKZBnuJWL/k/xwrfFajxlnpEmy/FA7yz
gSAubxCZwSiQNcowIv8hcdArrvdZBEdFk8W7/1Zz3Ms4ybANW/7XSnLcRMyAAsD4FfZLaYpmKk+p
oyR1Mi6wSHuECx4AuFwOHKEBi4jBrfbETlGE5tpLxNDNhWnekYKpk9LUPleUcEMyduH5sK0FV+w/
TEBXqVELJwEiCI4Y81j3eimgPZJ8Kc9p8liS8n3LD3zH6IIKSR5ft6rlm3CcN+GAYpUDTW3HILG3
izVx6umNttK0C9Yk7YyTKUvjjPJeGZk4eEiQOubukHJUt9335sIqexj0iN1zg/OG+bZwjica0pMX
7AYDfPaL3NAXmCvi+noGowUaioErzypqh9uGtKsbbc7TZDF1qlVpBmgcYeQHswZYQjEsQxOdd69r
FEeOjL2fjJnqGvlS+AiarQWm+t65Vv/ut1CVAEYDECTL1Sz663cIsXji4Ua6BaeFBsDZgRPutxlj
QBgrBU/5SI6+YQFvdQ7hQzrXwhK9fa8w4TUAS2eWnGZ/wXlzeUHudkO+RNN3/57EZQs6IeJRNdkK
t8Yc+9jEG0GvcwASJIX8+zQCux53mm/B/m1OU/UAenoq1FsHeU4b1LzEw1Bf3rOilpx/8SEDi4VG
QKEM+kvLivTWlGTAcpAgFD8qkjEdbdBx4r8BMy7GPGc4g/rAV/n6oEcapBPKj9/pHah0Ges478DP
9OpBtMA8hXfOHtkB9OdZMxfyq11tdzuZHLH1StSMgMzW1SqKg1AohjPafvjxGkCBh65aTaJ//nh3
DOeM8Kg2e5n5uZUrUci5boSQK7T39WGPhkvgpWObOn3JRrRNhFcNLWRml7+XgVAHIN5QOOUEhH3K
Xp5rQuYzTWy5SZXwqmK/qqE3/zUjPBaO3Unw/wqFA12bU2NHu8XRL6Bml7X7KrJM9JaX37p/avVQ
lTyy3bjEQBKc9XgzJHbrYD3vVgscXREofViGmdcaZv8IsCx04/5uF9krnS2pE/Hh403l3hVK8ESt
kIAj+IRZYshy9v3U05sjGgapYq2Iiz2psEx8DC6yHpJEpctpSlizR24LOgCAmX7zKZrekU9SyD43
A2XAQOROze8pqCPv3HU6Q1hNw6I0MSHRlreiFuQVKveixiFdenV6BMI1ZnWk51sugjOALgVbxd5O
hB/SF/9M9Q8QXJF0KSOG9YVuKO25lVdJ0d/WxscS7h3GIkTYXyLWdIKtIAwPljCktSZ/a0m60x0+
nbPsJIwEu8/rjZhUK3RFWDcyp/4aW1qeBK7JOIfTMR7q9Le2Fw47EMa7EXnZHHwcsr36+ozATQWW
/Eu1zGMxorOKZNg5k2yJURGxouxlSnXmhMuMRpKiJOVakxMYEyEnf1CsMOGLrA5Q3yhXDwfmPizD
Mvpw3CSphhcdITDOmzZIZBn/Nckwo9RPUREyetE0UtLQSETs6IP76nA3DK9IeDq2ic29vOQNIX8t
COBUFie5wCLyKgJ+KU0z21j2WZgWSbMZtlXpDkizOTJLZNzVqwbkXCs1R5H+pCJ3nagcU1GU5Zg0
u2Lxr2J/2UDidtZS+15j5cZugDPK2E5JBloKzWvnvYI6/+Naf6QBITacBgIBqbD6cD1BNcQ1POqG
PfzEQqCp09OlpXXI7xS/vsEK4ZuEEMhQXzFiXBUdwX1TjZ3OgPEzpv7pVR2x1OYVj4+7xrcdM5TZ
XCVCWnmlS3y3B26Y1yZbF6VZC4BGcz+1fz+SWPnEFNTGFFDbT2TqGhLKGxLuoiNo46WQcE+QgFT+
1LozR+l67um1veCluggpJuk/Jh6dGP+0Y2rPWSJWf+XZuHbSI6SxU2hZ6AqqVk4UFkkCvfWH8DHD
f0klTW9rKd0LfXYHsnf4ncLD7BOjHaFdjEEYOhVs3XAOxvJbU7h+GM8hf3eWAEb+Y8+P7x4h6pXw
r9gbFoA6A2OrT3zzc1itQsVooPhVLAzWOi2McYXja8/3M+6ZUD5izN/XGS3TvVO+rC/ktV0ulknO
9PvFsQ2TTcBzFoW1cWvR68DAbb79zPRJUrxMvzU/qkD3g6z9iJxqkqzoUlCKsH0qMmxqlfBmOTlg
mvjlWD7J1JzbDTf1+qJg6OXaQUNm8RRG9PI3zMnOvrspKyWFiUvMWw1dca3oPO8GtFWNQNvrEAGC
0bZY4q055VxODzC3jnlstpqZ8BtYvi9pcWmzCRCg2YBO+L9vRYsWoja4CHRSr+wKzgxglvz3cIpA
OCm3xRt/kDl0OcbImo8Oq7Tryj95WF1M3i0GORu86bw/MuIJ6bfyFo1r/633NTqeuS54Tzyh4Wu0
BGXjdsMVgfP4cvzgugWqJkObehdjmxMSP9Ea2iKCId8aeyb9SXnodNKVNxtW1wM11n+Qk4QKrXC7
97h0e40sHUctyiDDfWgSONmpnEgdHQdDpLZi9/j9JQmqi3bx4n1EipN8/Atc+/nE/ptlkduynOJ6
KMO+N67CZQub8zO+5w2Q3O6hERjt21RjqWVgp/aZUMgmp/ZRfSoDuN1P0T3VfTWnWOulAwdfYqQ1
9mun6CP88/ff4BfF6pmtxMg25vJIwVZNJkA/wkjIhuVv2vLqZUozMFtHm4Vp58b1JDIEE5jzU9Nb
YccyZe4AU5q3CcpSF6rxCqsYSbKWxOshoRrt2f3K7fXlddz1f7A1I/J/OU1I93Tk6jLPklwp12K6
G12NZP5FhZA5E1pHnbareKUO7760aWaio5PtGwEt/XoAhZakJM28X3sRkYe0XzyhAAj0EACxgGiq
fdch+9tpPxn/0EmBV7yOSPd/bTd3zStA89Cd7u/AzTNEcNnSaS0+aKDBnSeOkfXZFRsrB2DDRNtL
yeqoaZP4UpqK5WPy5UBHKFfLLrcsSjiVxh8lFd1WLPO2SbOfu0G3r3sH26e4IwRCdptSieAXpcka
7Tf8ttS3HjzsqTUnFKSEk8jouNk9gGZVnqLfxsY1uZmJ6ZEv3u17MoYtnOZwjqi0vpLylJhyQWA/
5HUNySNZzreYxHSBdEPFGVBtegEfnACpWN1ViZzjd+DhbFmwzrLQb2WT5uCmoB8EzfPxRow1SAbA
HlznhZF7ug3bniV/UTBaDiJjVcTVrPf6O1IwfWhUw2k09PLYBbx+htRzg6QXnMdUUy79X6GWy75/
Xv7N4/MSZeveh+6Ez3Ld2UmuxilEoPdWo0bfAo9+eEKgDahBTPfNOfS313iUEeXIa7qXwYWnMDaW
5f77dQTo6Ng7nDJU4Xgvxnp3T7iYu+HF96wEnJ+htJSmunRoVd45T8iaqLffA4kX1rQisYNqJEbH
xVSO0hrMPoYCDv7xYAVDjsJamAmPhWJWfGKaFzJydoSJhPnWj8kExEuCFljTACGEDbP4OqNs6h4t
WjiuLOZSr2u6eyt/9pLFTmqBkXu7uYTnmEpD8hUXyb0Ewa6pwud9oFeUaJEKNy1LDZN/SS+cGx8K
UGT4lTV+QBEPxt/1DOywZCb1NJXCjyP849M0EWNCBdjfG6HTHdOnmrwdpj4hwjljXnUliveC4q07
609zh0NOv6uHR4us2gnLHl5JV9bqRmQQMsJxtZLlSdOdL+jQCqtWScnN+akOwc5Ea6FzaUzmBapE
wFiE0f83SvuJnG1pxGP07wsBEOtgGJRKI9P7lj26kEgUjvuEHxbVO4oWaKGpShDfN2sIuM32ndYk
jyAW51YGwzUWmCvIJFsJRjkEUxeKZvKS0epaYTk40sT4wneLX42gnrJP9rLsZ3FGn/pMAmtQjAjV
TaYjAQDH2BaJ4q0nx4+HRAhpOXwMxvomEBXL7/IR8iBtUCXa7pIMRL8y8VoyBR8Cf71HwPpaOSmQ
iXdmHtG102hfROXYsK+6PG+8ghen8EmqEK4Y5tJnEFwYRFWixiyMTOjYSI4U4xLgs0/Ehg/8wzF4
Z2YxbwZX8aAjJtckxy5p2Tf4lrxuG4vJmsIULZSJvd+Ww2tDJbvbAtORTPXL6JGFMfaMtIHNE1dZ
8Ly1BsAt9uce/JTEBobrX0QhwgPdLsepMbpYuArA5tHxlUlIhCgo3+SrHjPLpFuxj/uVDa+fy9+4
BySD0WgHjF1TMRxi0H5TTrT13iUcKWZzxlOd4spy3iLriR5SLJwBiusWbPshI8g5eCz2AZRmuhkT
JA7TKujXY2eViTWP4t1dx6iYxgVe9qZHk67mX/2C+MGLIK1lZlQSjEIaoLAeljSN94CpUsZe2wr4
cO8908Ay60U9DRO+k8jYVB/6goABP54vKB9zmFWWbgF47IlK1IomPc2kzPXBgxIoDcrZcKJnRO9T
ohhgbg09QBbaS/dNhnw3zaOK7Z9sYwUiDTWQU2AGd8qmapjJrkjX6fXbbflRkORsULYo05Q7NVkl
g5dtxR+uHaljATX8o25iyQU+CeTUZlCL/hBvSTRf2i4w41YgoYL0+XuTucXKpvU1cEMreNTSdVg/
9PP1onLnAJ3HkDuPk8FSEX75rqTZr+EkG4mIJdFkkbtM4cDxHxyh5hVIgS3tXZzaVX7h6MiQ6Wdu
7+hv1cvu+kJho7bl5IaYLu6y7IkXnBSgFOfMoct30ZWWaE5WgrezUV6coXwPLjDO8bcpYxLl/5w/
G7tC7eZdn7YOmNvVB/VgEzQLMVG2ZhF2EmQsKUIqCWnkea95f+TUiMs2OlNXxYdaoyMwqcemNbtL
TBbGMq6untHnqMs4qcxkLsgeo46uIvXx5STiwWT6u/Cjt6lswtGhhkktcnTYLCab34a/j1NZhnoZ
mRZfL/ZebscgkaLJKanPUABRZIjQDGyaChppaWqElGyV1DxYhO7riLjm+1B1YXOVxf3F37BLJjnX
RGP8IAQq+/+Ux7tXzJIgWD3+T4BqVkvawJs8JDGEfWdx0mNuFnIalw1gGYuJpEfN/tRLmg/DKCgM
8WfPTml4oF0zBdUrsJhQuv2zfZXOK+JEJ6a8rA9QWQhHhYp8715B6Sze57SUL9tUmlEKDJv/gtb+
hOLOMJBh6GFE6KTpyDttHG7CgpO1Nk8M/FxHrL4j/MnnjOj9HaQ7F6n/69QIa7njh60thk8LM7FS
MbBm3FeKVdH5+Z8l7U9llfXf8lRFD0xOC4OOo1+6jFDOGkxV06IoGsm8Tt+paul9HE3mTAYXM+lG
JsykShpCsiH3kKqPuvS8FjWgwxnJESZTShkPrdTTrNbI7UnbZJO7lq1kfxbUplcjbMHRTfDEits1
+1d/OPPGc3wqnCjZ/qI4wqZ7mANCqRal1liomiXYd1ObV+oA1dydo9F3c7xcVpth8+Z43vY4WvNY
e0VKGgDfKbBmvoaItw36GppFEGohbTAeIjBMQAQQDmUY9kaGkrFi7O5NjE5jiG4mwp4kfYetET0I
25LJ3zveWQKXLJEPNhiY3z7xV7buQ0HFFoMmTsaeFT3pGCHiNpL4sbyf0YfhnfzjM90Xnq/FdKyR
B448CQwBuRA52LG1QOHqDL+dlBL4mQtaXqlQ0zAlt1WXDX/z+w4Z6+YK3f0jjK7qhXHmgzj26zmi
4FdlToiZi5iceRkwyGoEzICLpewWAl3mFja3y2JfAX9rd/4TrGNuQRJ9RtucqCypKlxB9DyqbsX6
eMmcHM2u2y0JtN2yFnKae0nUep02Zu7FSyxy2Gm0LHXct4TcG4rvgDK4UqWVyjAvlz4T0pCgy4/T
McVbXBYihsMQqc15bViUJTsEj5NCpSspjtOUFIzbpO9ztuBejbypz830WEj6Kl2p1uqnvs1L8N65
4NViuEVl70QRQfjN8qj7q9l7bAMFd7TjtEsBmdrCnSHdh3YBNykRETCJQFVxtJd9ICqha/AHjIGy
0OrPVpQ+HCjeur2QwfoqZlqQPDRFvpALNuli+P2laoD4wcYPGzOjVDVcEf1h0HBao6xkLcXgcMx1
wHrP8XSnEdofCwIuI/TD+KtPSnHO7RU+/yFJ5kRzjbZUdCr34fYg2df/Y2uPNq8MNLMWuyXQKekq
PZRKSktZGJ3Q38aV+m7mEP4g8fNRPmepPKt+w9rq1gLRKgzMYNHDdnlCFJNtBBTYJM1qs+jLlx7Z
7+fXGY6D/nwe/LfUl8CxYv1DRglYSJln1YAwCVAe9znfZ+pNbJtEcIf2qyHm6dGeE50UKo8bbHLy
X55Ma0gdaI5zrVRoF8aKAwlpHLCwgHHNcFOjaIhpiY1pRr6S1mXBmOpmaPKdn1r+lzNJRl0WJ4I5
OvsdYJyz14YW22DzRBZa1EmCDLJC26ru9BfaIprPnwWSpbpLsRbuql5m4jNWEpUS2QCL16BCFNqW
jAahvZeb9DOO27nUlJrIydxXMTcpzqvi2gIwWhOpph9WQDfzsv3qzMMFdcnCPLD02qZXY+d0h7HS
dhdbErRL4Cah7o+Vk1ZgTBWge+/CYJLsNflKPmJcpwAFwg0i9iTQn80nJ2miHSZQ5P2+KtBohNtu
Vo8Hzv8OJUeGhWVGOXPl/rzExAz/PGu9pw6UQxVTbR/WVnx4KEwpoRY4k6vXMTnnvfIgEZuKEeNh
HLESp17GriCXVj1mpMgvsrxrU9Ys9a3UpEWkJbIOI52QqLTWrq+m41UTynelpnP9t6YrvnP0eg57
2o3rMRx0eylRkts2sMm2m8zZYAcyoXCilcmpazvLgcR62OU3j+fdi052JVW7DFv2zP9pT6eceCk2
twnfc5CN1EecIg2L/MUV6QBmoKHLZo7L/XqdJ+kQa5GctrT7BXdhhUmnTo2nIDgUMsH4tFPyvRjj
p0AVYpFWn7jVsnQtL9HIShQ6m3Vmhargrm+n+RgusWMC7XCSactsUYE+0LWPtR9aLGTst4rs3g4C
86Si11CogD3dkEXT1frR9Z6uZFWyY8+wDt+pKICfQk/e9+XuXcu66LznI95GY/rjPKiaSpwiHCZ2
mJtEQpciBXWrjQY6dWL9aQjM+XH6JPfynSJLXoXECY1xTcdZ+cg8XOraPCCUg1kLdKmDe4eWvfj9
W4SWgrUelfjW24/D1d2DwW3Th4LrozSOFfT+EwF5kTzjffZ1YnUX8wREgLStaIWRsaWjG7TihMQB
7wo8RVKHj+1XS5kid0IddW5/kZ4l1wNHjNPisICkASew6Ot2KsonV16/0Qitky+dc3EzX+NoD7ZN
x994+SdW4yPcTe8tcOEv189wU2EkcRya58Zuf2SrYgMhEi0VVhQAmEYUfwcVKH2/6mARCqaLMvvY
jHxb+axyAnOKoWqECN0k/UcFM4MJYrIVnAXfWlA0fH+MQjxp1AofUe5E728kZVDlBEdRhRgez5gk
T2q+YMq7VSMb3pToPjWcPnhrTJ8pT1RrzQoASD/7xpaZeZ+AMapOQhhK5bxlaa+xL7oVq0xWBJlW
vGi26a0pUZWgHZX+S+fXLIl5kNyr/OC5E4ElAif7mqfsUPIyqz2b6qE+hcyh3JZ6WHrodTv+CvpC
6+WHXAF3dzAK3D7qYhewTzesxXulB27Sm3OxTrsx3pprokjXk8cv7/WqRwITPms7FsvAcOv0rTwb
KK73WQzOiJE3IY1ery2btBJJFTpgyzoi2tuB6Ioq1b//mhunozRFuIW3QKJ9iT3tZM+pI9N1aU/O
krLvsrDSpNCVeta0/0/72l/y5iPnpuPEKot2SiHgPHthqNw1aUtvpOMC//mRpUSKKyeGhSRRnv+T
KkNltT89tJUTlhkR7Y8z+AHyHhcxJGqwxcmbPZsFb4y495DKRrcV03JoKVeNgN0enNbzITvwwrOW
LLWyA6bg8URB8f50+e31dOJSZXRxC5Ao2SfQInPQ+bkdN0D4r5NzWDxLsGbqeocxOpd+WzW6M0wn
x0RRnTWPfX4hOQsYhnSOIjaXL3sS+N17UEa2fEHyo79H3x7XCXeP+KgrCJPJVMh6cKmy3gSUfA2N
uMmrmxemRUFzveHiQ1xR6MeCyBs9wW9iGWN6RZsMQI/UMTr/BzFebjieq5TdSu0GYNtsYy5bmehj
Qq360v0dx64Cz5X1WYF3IEEqF+tvCQOcT4nJyGvjHPkMGXP9aDj1/H4tArajJkzsFS7hzyR7u1QW
/hqiLRJrTZKsHs5KR+TTB193uOJ8vP+/qVbmEmDEvpqQUXX1VivJDGWNaKqECgkVM2pkJ27K189A
qerNM0FLREjMSoOu8lHk9ybFx0qCyjrsqDoQNPvRvud0+DclYQ2RB94qvFszM4GfKYFAuhOQ/gxM
daV0xz1UVn7YDmMO6aUfhhdSAet50QTm7AFdnYhtgkcwiXmP1dElRbxpnQb5K18c3yQvOM9N04fG
sEQPAJyuycR2WqOJI8FEgQl962oZWqDPphq+cuzj3zcC84+7FlfHc3WCR0CsaAfVTRib9/Me+UMj
zlSisbtFZqHhvsLVnd1QLQZelY+VWwVXRGmJ7ajJi9zlnoHxc6QTbIpNyg4SDjckHGFmnpCtuNb1
jrTmSmVIxBsYkmtwxtMRF1/7AvfqIjmQBz3bc1r0H41rZ/VEhOv/8BUy69UVgb1QLbyZ9FDHrxTJ
7Hw96GXMAW7dWgAQ0VAxsmkY6Wl2Hbr9/KB6klgDhLBNzXt3aajU35w6ZnK/ARAnlQJ7bg5gH926
S1Kwwq7GGZuYBAYc10lx2e2zIOX5VV19RCcq5SRCZQnAtonVeR8di4B1SwWsE3D7I6NSRiixv16E
a2QIr+w79ZMF3RhcJ/WLQ8fO2xd/HwF68GMlb1wSJqpzgUpXOkHvVo/Ek1IcX+ZYHbtLXfekZesy
N+l+HN+/4OBYoMSyNX1+wbMuSgo6TS/tqaFITywaN2TKOB9XnRiZPseJFtp2w736qBXp5XrLWhx+
k/IoysKw/IqsIT5RC51x5gcPSPzoDrwCtyftjk5+N0loStASGPFb7ddDe9nA08mNhNT5v0DLvmKj
FXROTXlTIDJjqJtGilM3C4tWone2wkXlKYoRiiXsnnaRaYadD/3crj3xiVr3c2YSC4U/5udPM3ed
pQmeamVJb9xH/jOXrVZ9PHvUeCqFEF1cPx50chmzIrh69UWgvamSQBm5nw0BKTsolgMwrZLAxo5z
XK7kakkH1TkLkpY/n3LVROSxOSIn05ENKAz8vSPSgP8qdoCsvNLtFy/HCUbOhVCQSHX8avvIY0KC
SB9srg4ojgICnEhGu5EqdCCkaShfs9r+2/cZvGumnelWo+1BGT9XMa+hIszgdp9jdfln/w6x+5co
NfjtDjBDpe/e/idcSCcJ1+5MZ5GYYmeIRIjsNR2tPKp9za22a6NnF31loW+OlUaM0p3IXaQfrmhj
HPPWvSt7gldCLh9AqRKNKX2DhOb93Omfs0BOP2IhzB1uwHPHnAlnwzbTIdMqqd296GUUA24dN4ba
G/BNJHrd8e9IMsgihRCgZvF46PecewN78RfxCOeLJd0RFr2Gyff1SYN74ZLN8rV2Qsu5IpabYXeS
xSJj7uRSJA3CL7TIHk/6Y4b9FEmqm4GjQmxRXVVpJ6AK3pzDF98N3y0U0WU/+mQTlTzEv2Xxck4n
tc4S5lN/aUjUxIBnU8t7QdwAuofhnD7tjk+VIHpJPSVONHgoHsCX8tUkrR1YshQ9YiPyEbfdBjlW
Jiid73izf31oMrGE0b+8sTsGGkS8oLW2mes9lUs9XX5m9wDUCojhqVo4+PD04QqZJyqKoIkDQ/Ho
3Obb/Us/CZlZob8csH/HKDXyaZE39fvhHW9EcgwW42ge+M7ED02XGDGKbNpblbcyQ5Ipkn9wrG2Q
OHXSHHNvUT+Aal9byXLnG1luFNVMwAK9S/PV0avDTE04+yL7t3z1HgnB8x1kFlZ3f+0+Xec0Exir
0WWpdWC5X0czDuS0mdwHPuyZk3FQgnikE2NKWnk3EZHuJLx8oj7CsykpJH6FtzQVrETOapTRmY98
pjFvyF0idT22YOzCsQKgYZ04geOtI4wOOqQzJ/1DhKFu8Qh8PlOktxYYRcnYby9DbcGpWijWDVqj
upUFx6LEUndaRFQ8sq65uE3i0y9CNJSMy+V1uZKgiXCQxK9b3/B5BwtvKkuhYvuUaLg593pVUDLs
INqY0D7sZMLKhk88W1n7aVolsNmRie2i9ckB80bjGrNuQxAAgyzsijL/xALvnGVPxRYuoJ2Tzufx
755qCOuTzIdLRoMyl8oUA27lXjcdAhYbEs1f3rUt1zMhYPRkCLtW3V1pQWENlPIQa9TFRc0VJX8a
BqjiZmzXmdiLWPIuN79k8ZKFkigvjBRbRqoGXz2ivsc6b0LddLtZdHb06mynvFUyge0towyGoW6z
cQA6ystpS5wxUmqdcFHKRuGBm/bbn7toBKecxIC6tSJPkyjY0k+6luXbZeNztiVq9MWRJlanVrNF
5lhlTEtcfalhYcrMyZbnPSr9MLdUhIfNJbrgY+Q33j6/xAzlW4uP3hG8UCXDSo1lmKPYshx5EP/G
D3FKTj1I+y0Ki4FstTbOvoXVd42abXbVoFmWX5Xc7lu2RTQlR42Ze54osKq2ykhFLqghFUQT1OUB
2ldiyqUZu+2Wqm1BhUI35cs8/9wKIoiwLmLY1V2MaaS9+wQ+BQAxaZLvZyBTKyht5YiNtQxqQj0i
2yMIMOvIOorp3/Ls2+ohEfvOBm5QjhNQ9VYWCko7cnLgGGRjjus2RQf9K4S/l5lkpba+ogqN0BQU
2EIxNVx6PU4Wd4REoXF5/QY1S8Lmj0nr6Lp+jYwjnXq5a5zRvMfIRgVlunwm8oDMpMjPAUmkYvqp
KRdD4qtNj/trgb4WN5nCRhZz9/E87P/h41s/q9ZTrBmkQiKNnn1NFSx4MWFB7DSpE17hQFWMO1yd
BkhCauKuwDMX6W7RHy7snekWbtdYjuXNRBJkKBXMJNCqq4La866hd3gLXKXu2XlXg/nLXJOv5XS7
jr+KWaGWsttZKkthPeaRkeHjV9lqc79sS1eH7sK32YX6wADsFJeaF+KVr/PiHa0zqO8oYokWAxaq
fi9OpgIa6yM/6HuIzOM6SMH5YacSRvmumMeempqoCgaODpe7OwQXJ8letcgmfso/IHG2mifmtzNT
jFTzymca0aPx8UT6OZn3YWyjI0CtBLaoyg8fMcDFgaZmVmcEruWS8tNESdwCzaBVgPX0Yhmj7GBX
G7DVa5eyXsjXCTy4TzeLHzPKJq8HTu3QL51tN2FKkwHT11DhEobLw2RaQP3QdcqOrB20bcg7nvwH
UwR+nCXYXxqg8JrtDA6pNsJoU4mUWHNUD0RnduQkcMR8eUORSwz+JvO9yrfYjQxdc9J8Hr08FBAY
GpD9GYtpBEebBHLhAQkrcie4lw7amGQHNTLMIAek8pT89HGqOWeAxE+1BJvghMcf0/LHDoAvD3SO
I/HV0aFydgyb3RsPg+ZtQOu8Eoq0Wb5Emd3o6/AKmhVu65s+VDRO00ygSAmV7Pei5Qz5oDCkqWg6
7fZYCJkLujg9dVl9H3LA2zo8ouyp2+ENApM8mGfrUJxDyGtmrWWGMrJ0JzY7GusqC7QTSybUaVmG
WNxZBMG4utLi+bRSi+Abrtpk0gIZavhIlkuPOvQsa230ftM4ev8mard1yg33e9RZdxopv0mqTW47
n4rl2O0MN3ZqDjsPbT5IATgqg+5rmgFbHhl5VxNJjaqQbKOhVo0OZIW1fXYjtxDMR9kqtx8e2JD6
kMAaO1ktU0lFEug7wDHlFte/UKCvrr3Y375b95K/Y2hWi3Z3qf3hrYreZncRcNVjzS7tYscr/z0X
T3M2xH3dBZfpyCG5eMLVKy9dS6iOpqm1UT1obl5vVrMSmcJ/PJQZYVKESc7lbncFPt3TknSEoJ/K
4jGMb0gDdV9BQbHJkMYc7Ln/xgN0HuwrNPREyPnVckEczPtPav7PZoCnH4HchZLnzjlqO2WVbJ8G
gAbUzjP29V1XJByf9bM1rEdSFS6CdWfe0C8OaFv9rh1ngHu33ukjCsihC8LS98/XXBt06Bb+ItyG
wQJTvC33YSgcS78ATMMZpvc9j1laaER+wYEOh74Vitd1928EPmYI3GW1ODMRbS8BGeM78DMJQwxO
KIea0yCh68vTLB82i5P+hr4euqbEN5tK1J3KbbrLS+imnKN7g3AnlUs697jmTLePwmMHqH1pcbXV
6GhE4Lns9DxjFvNkmd8gC9qFIymkBpC4i5KpZZ1066Mj6n5Ou5J6d5fFQ7TLvouhWyWXBCnSiDKq
15wiEcaPASNegDRqdF4Rh9yfN8uyA0FNz7k7+7DHQY6GBgf8+K2TbOngfzJbBUn/g1tqI6pNIczF
WjWgJThtndqRtT3I7LTCKIunxd52do+GpQksGAbQLbqVzxwyZp+KlmzaU4PAR1scJajLq4KWQUpB
7c5y2hRuQa5709kGgkAdL9AMZYNALlbFb8eZnxTfG2IyxZpGE6ADVTEYnKIr4CaOFNC3nG3I/n/E
2tAnryf335V7WsHk+CtVjk1lx9Ss3YKamnZRaNNOs8QQAdueC410zTI97jEuPH36hJwshWX4eF7j
0G980x+/GryIMFCsgdNbx4oTAXMnUJrDLzrM3uSxKo7ozojSwsTIdjI71PykvaGtlO5b4EkSDJQX
Q9Kf+yn/ijjEIEjvFEyDYmHeD2py+/bYPtzuZq54I/Bq8PlyCLDUqHjb5F9wa2u5/peMaehkOOVP
4foe60orbZWkkXu2nf/tiUKYS2ojr4UlLSjqBHWuavYD15YclO7e3CPwE/q+1CkwvZKluBL+jQcN
q7fdRvsWj7o0siOt8+h98v8Q1LG7lCsx4vHq2pwB49m5ENtUlX+iv8A1ihwG6KeDOjoZM8eMor5f
cQPYxZLa6phirDYaZ5EQTBOVcl33vLG5zf+ZJANIjJ6AYl8fEGbfM0aHYoXRQ1rBvjiboj66kgWx
DMvw60KNC9YNQW/tMojyfOqfLgFjKCWIePnbctQgz8yew97pe0DyqL5MYWV8YLfYdG0zJbGr8qqv
DMmlxWG67FwO6poqI/9R8+s/B+b9g7WMMigbjOIbJUtAgQBEYNwUQrJNKNnrBeRtxy/ZQSPOTk2i
8k0p6/8kpbC/GnhlhrbDu1Iwgi/K2Wu2wEtIApg2RHfzXqKndpYTXAN5jSEcqNryIJF6HyFVaCx7
rIOTQxxT6MzPlc41LVXxUyUQ37IxgAbW8pLpf8/pm1UzX0gbQ28tXy7nyEZZGt2JJVEihLbopy9x
rjPdrzAY0buTclX3c/Gn5q9NghVYFjPqD/YsXviNweyf6k1V2K9Lo3f8rdXxBZN3Q0O676TY3vWa
KzBbsf8fxfYF3uIg4GVgVn1sVsejDCzzVd/rHpOk18xk8x81EMmNuubfORAcGipM+t5n7cb3eNft
z6xakM96Xsk+xlB1wS/2pnev5A0dKWnGDgyE7cz7bJOTN7Zvb2ZPvgEVcMskhzXKWYVnaVJqrEqA
WZSNmLXe2xQvw9r389skkG1FF5f7KZZLiE19RK7SxA6tuo64fS7tlpv4X6qKqB9MgFv4WytiCfzw
Mj9tfDIKP7Xfa2LJGibVfNu2hSOiYqI7a2UN8pdSjKPX7YhMvSfI7qQVodEwLdBudVlDWrMxOJJI
yk4gKN6RS2fxz/lX4i9kws7KDvGab3I1lqLl0KcesAOjETBvwlGZwlTrye11GF8yA+YhxSzKeYIz
5pyCCnWIL3NM2uRZlEwGZ5OJolru/3usgx4jhqQB+DgVljLPyfHKupWdjtuCxdtHOVJ7Ay25XIL9
J+bmyUIGWhuyOAIqCA79e1BhC1mgDQOcDxpM76B7sTzDUpAGcp+LGX5IUjHgNwvsx1iQgROQ85rs
kxpqFMKaRwQiQ3VFLiAAmEsDYsUP3rRh9h3pqzEySQdCIUuFwuS0jRcCPmop6iYuPi4mMNmoMnIS
dA52w8nuM2QfxhTR8WkOBBHpLws8C4RVw4Uc5jgKUKqstw4lQir95PXd9hHoRo0monJ6ZoW47ac2
mVD9hsjvqiYrY2+Jq/NOW7lKvlhw9jX48ZGN7TTcQpFBcp4hWWNmPzMsYRdHvIGuNLL6Yy/JZtSm
9mBetzj9qVUcP/s8/VmSs1/MDBz/fM9qDYjlc3flD4o3BT2r9j+N3syoIX8uBp+BQQ0uijRitMij
iUtGmUUiJudC1wUFpLeH5lFuUh3mcEkeTJ6oGc24CEyve6pOrUtjrUAcpmUm2viFcA9ikNJtriGj
PiAga81zScaP2M1OYwXkot38kYPQanWGMc+tiGmUkXeH4/d7SfCwd6EBf+xZp/D9/n38hGHaArCp
kxafMpgv0A6DPGJgvlmrn8AIv4bOU4Vjv4dcMPAES5zVZSJ1SQ1v4VNvRM5x7RG5G2nISDMe22AZ
0B36YXoEeXGBbFkdhy7kE8e9zkDWcbR9AA5Oga72KvadoayjVQdhT0A+anwXzI6GdiMIplwiPTAe
YgRRrwmRjLXGVkVBxqzPa/5jw+RlF1vdgeVYGpnYwIrRgcjdjhsloNln/954mB0vv6+wfxUYUXfR
jkUZyBiC0r7TA8Pbv7qUwoqRFylbY93eTNkpG4s+9Z1LdKU9ULVQQJn8lVtOqO15wB1q5kGx9PWu
ksKRQ6zyKxYMl+Prr+4lOvdZHl2CWlQKJTgVKQsKQNA07+N8jg6tud4aPgMuMx76jWCGE8oJcJdA
Idxcllqx4OdKVOanH+Y8YEUgoeVQk6CeOr/gOC+J/syZZaEykdw920RDF7ypxZxbauMUbIcE43sd
SGmHc0T0fcJTl7I7vwjiSasN0lpf6Al/rn1sXSVa6ubrTvSfN5E8DrzsYlKM9RnKMe5/4sxfa/Ha
XhFsqpAK8VhKMNuvSvibpjY+W/QKVp9q9WHTHp5UlHsCB2CoY4O3i1MmqeSAn9PGyc/fw6uLn3j3
UFRPGMhCWKlzF5gYhhnoPq+gvvnKVC2lAj68l3Fknu8Smph4vTf01WpjUhlmjyd4q924peGTIg/n
v7agyirqVsZt+6ncRKZr0ld9a5g95GN+kaKk9tSqyYrqOSxBeFDlV6F6zdiJt5ZozsxMFuKoQTNf
6tnuaCUfFqgL8qVmUmk5c7NSHQp8HJQa0XQ+mKhmnWnox5eTBwXPeiwVBUvfKEsGQ2NAAk3+jnj2
mJCYGQ+cywRCJ0pbDqJi6xBNwEctzZyEhTLRrOZjOYupF8YDmIQ85o7Y0wjF6hWom3wCFpn7XgCy
GWXGSuuWTUTN5A8EqFp2nRMgK8vwuB8/V4+bifcMQW8WkE1bOKTu4be8ZdnDwchv7WVD2C4BZl0F
zC8ta3ReoPgOF3vBDqUeLAp0RGZhmol/1bhLu44ykUcmmaSz859juAHeCZIajrQ/v2E9sfiSHCbZ
+M4foRAedbPmSyLCzVfxICuPv1TKq3ogjBeLqxInFsbzBFW8HuWO9q3KLvlZahxPL3h9lxkRX/A5
bMmVZS/KENwhBJ7sIdWrwp3gj8Y/u5DKv1AgJ/Hd4eeoJV9WePAT+i9O288UsyTjifSKkoV44S/B
CrG48Soc9uekSGenfxo/2NAY6z2SFs3wiTMiGvQSgy3aMfTpFk6pZHc/vaoxUOCthwxfkhlyMtyr
LY5P5RlsMNfDorCvj+R6NqYluSRqb7sdoU68bX+J+Qj6crGeSgpd+OwMxA/DnrcfpPzbENaiSiLK
h+36SiSgdvNuz0vOB8Y0SXa15j3EQAhw4QVcoORNZ5HzNmAeLl52/8HYgeV1zsZY65eQtt7sMii+
VpRo8/7RvddNQX6doNZa6fO/QmPxc3SQDJ4RvY1LCH/EsDMw31r814YKT4fptzNaOZQVOzBOreHg
HwpFJhJ7WnJeCLaYSL5M/nJe9vIFIx2ZDBzhrr2fZBXp6t8mio5/f/lVuMNVC90yskT5TxixhCYh
R5lmMFethstiAmK5wmSdSAIwAC4gUf1puKX/7gPilZDRp3ufeXX5bZu+ja6bnwK9xbzFW29RmFub
Cu2QwTLIdgGcFizO1Xar0GL20tEFY8CEOGlppnw682d22M7vgUuAcsQNgCVBcL1gBE/a9UYz2Uez
bBSD825zZO4GxBQnror7CYpRmunff9MPHnHcq6QBtkRS05y451BbLT/WcCBOC+pcg/FAvfjmK5aO
NgZPn0623En42uMa7IQHdS4JU4RqPKdrMXa/qj2nROfDloZ6wroowdwEqVGAKhbNQ3IDycXDIh1y
U0DxbCKrxK/VMpAJ2a+Z9CLFBxDYmngb92pzjtzL2pCSkcDjXOJ85PYH2PLRtOq5mQ6PfvqpIF2x
P/zVd+nOLk02OPCTQZxrYstzQ//VnZSrztxap+2zSwGlo3PIldcGlhwcV1mbShEYyaR5NVVMn39B
T5Mosg/TRaC9AtdBnxBhHQwV7M+OjRQF85THFTCy+eS8o36dxmZETirGBbAoVFGGQaVbZDoreLqa
mgK+e/rd+fVLCrauUWaMwXjDTAwE+ZDS8Bn1dfXROY/BvFEVWfLFFTUv+dLOOXI3l0FOVGIshGxm
L60Md94oO4+TRSelZMdLulaf9+NctFTbVzBennYjc/l0aGtaLtb/tl+6x0s4CKkd2bwa+PnsB+lv
EYPzpWwdKrWbRPyBSZwEkgyfY0I04lI258CyMn5DShwP8g3NoUMlWFN1Niqi+bGHjUMluUjNJoUm
XW/j7/rnbjpwjPZYTVWSqGfEctLqpjcm+1E5vkU3gk/GFYhu85HhcGaofGjLbxphW2QnbHqyv8la
/nAABWw5OF13TR2N2fCVynD8qzgNz2nuw7ZuoyCO6+lckoHyOYJ/aSLYnwN/Yr5RauItluh36v9D
Nr7VDyQ+CZnxE3ZQYPlvINP02MCbclb50FxOng1s1aHY1qZFEilhFVgM0C/XP4KEjtcMdgGHsPqx
66SktDqQyM7NSSiJoATOc/EIwV7Jk4xo76P28LMam9ibjdmEnaKKMx9PLJ+bZ1kjdUYXMAcERBxs
ae1VAzPUCel81+okBvXGEk2G4QDOAanKT+4DG+8MNJO+b5l66koYwUUkbpdvIk8GqcZtFw2ISVom
dtWWV80O0pbSX4vqB65rHAtwHxycn+8EX+spUpGRqV+xtjlvCs4U3d5J/FWnKEBzzglLs7ER7IFB
eL4ye1+rqTIIl2TEHITiC+KfO9SN/Pbwa8DNuqc3WXlrxfwhZLLr+dgIk6VmYE/gHpiReS8siV+x
oJy2kvoWlPYjOnV4vK10FHJvFUDFqzqDX04pVzavKFq/t3A9YO2TcgiOUnTtMOV2nvTcqkZDS7Lk
PVWtjiyZCRKnS6eQYEEL8nIsF/vI1Fd2+ZSeZiy4nJEQBTK+Nm6kaLfz62D5y8ZN4ROsADURm2MB
d5im+Eex/S8PBFVcfA1xgqzL/CWjTCdf0+ukCQ+NkwAxbMFdKDdw6uh3VM7LxioCZ9ATT2vAMAEk
N6x2b+6ceGt0gYeOeXUV1JuaEjA3kPVueOjoMpujX9vtXZD/38epeXDQHne+BGTBOOwsl6w3czq9
abfo48VDOYIOu2O387abZG7gKaioTcudKuL6kuw3a8gIaO5ZgAzTu6DDT3v47c3gXpNvW2Kx1lOY
6zCOARjikBPGbIbeWMdQKNIGRf5wrJtiXTQHrwOCzsmEozsahku1C190G1j88S9+9JkJ5Y3ucVwv
Fw/s/wt9hjvGaE9t+nHZ2gs32SXlIKKGPACf0N0o7cr/x8YLaEypN/eMLOqbFQk2fo12mXjzV3xN
4vpx0+bfaoSK0ci72Cc/FcRzt/30cCqZvm9KIOsvETuY6fkQtgybe+b4jAnXsVPAqqQxD91QN/Cl
aM6ZAOu1K3gqFEh+gie05v4Rn2pwuJpF4EvQ3Q68oPpxnN4wJSWmxZ9ojljYKXNpuUlxyWFUbWuV
Jg1Kupfd4ZYUvxpVGZinUSde/nPPFQyb7KmSBvrCB9h/xEMAcHwb0HliRWLwVCF6ECCSu0SBdSsx
Y6+MlaSgw1bcK0BhgvQqg+TWMnG61U2MaQCth2L0A/gi003P6mM8vFxwRwA1ITir66eTtaLuGPZk
z4d7EYgRVhe+ru5D7C5ebPnV5VNoFuGJGze7+v5AwTm1T25SUU+DqPKpU0LT2xNmGziV0XopS1pV
U7qdX7JedxJUcLgQPpHL3VXp5G/GO2YUtcJW8l88ns9Y08xW1YXEkwNJwmR9xXvZi8dghuZCWBDq
N0z4VioGHgrKpHT8gwV6R4mh1nUG3w3sklEMgZ/7YxObCPl35mFESvEoPCYBSVoJk3F3VcVBlkFh
a5BTfx9JdxQs0Cn3yNRmu2R9zZ6q+yVpd/ToDp8L55CbY6XV9Il4L7zHbA0TrrHYUzbKqgVjawtF
amat78aC98iHr8aWMn0W0JmoDhY940jyGY0HW0EUfsQ7fwJERvQMbx2w2j5dmof5uKUYR5euF8hR
eFWEF7QhCLOspyblVR3mVuWzyi4f+o6crB65me2xhwNYat4lfwLAHGr57zPYofUTrZRGHD5I8Cdt
zngSZMfqm1WCRmyZcJSPIBW2E1PoVXcOkq5PdAlIr1XXiNb8wPaFiLoysAm4wF1F42YHK+P5KkW0
GSSIXKx0RUwDzS5ZUKfvX1ya4qFCqJcNRHf7YVB97OPyFdEJfevgg9kac6k0uyVaLegtxRTsIqJf
sQ3CbH2EEiZZvNe4MzFo9L/WTFWIlUOEMuRjyOh9lc8gUmCr5DReDyU9ThZAhhEICP5QeHeH8dMP
HvjLJ1Qvyat1JKnWfhD2qQRQiu9lZb9pNKXJsxjwOAzsUJ0nWe0rlAkhYNirrD//N2snzdqldw5W
5OeJQdFReO6VHCbKv+q3kPXevr+Ma8p4jitCLvH3UAa/7yA/D3CwK+gtjudb2sK7Xk+JxX+Si5AD
WZV9E3auOhDsSXKhSmvWuhl4meYRbS8UyfhdzkwN/Px+oyIrionheWDRZxDAkSEkdTtwmI3QeI65
6gx2G7G5lrTdLSNjxMnpvsx0sGBuVB/H7veVxoTDg6SUwHXlrNtFP8bDRF/sT069Oc76S0XK2q0Y
sOKM49KSU1X5zDOdSGZzAnsCG8NC6a1lo3wZR1TaxnwejVdgrD96S2dZCRa+6PxpGFTCIqNYN53f
iS2N55/AnduV7dBhezdecR+X5ZXne9AjVKp+5YiMzkjEeLVdZbLW5ed0YbcJ9qBWBpiSEA2JCSgR
cm9LZOUfAruhvYtpO3WyR4E4FPDDWBErcO/8m1FtbHjKXaxIze+qSBDE9kx8CnAowi5UDoQghB1u
MucvyziF2O2lw3wMFkSxjjXHL9Z8Dv8yWfYU6IvkHZrzVYgZw34kp8rRAgm+W7+S2qxDvSFLUeqW
JLlqzXHls2pIn/ICNYmzosgV3FePOCZNMNu9cUwo/KYqij8aLtK634z0c8XncZ4XK6lGai/yVc/S
avlVZKUMMuKGDeZCG+U5czzBD6G/wP+GkJOjM/SlezV1qGMfyTRv43hdm1b3x8lg6MMM6wji5SDj
6hjMP/8wbK7iIxFpK54AJ4rINsaokAdohOxVQM26+Na4h3f1yZ0BuDdP2aP+BESkQMzdPJAmrDAw
XVj1WWt2p7QjQpthw0r1NGfoB8LD27eLn3NUQWCNpVeQaqGF2pwr07PViokxyYM9E5EzYG0CIGo7
Yea5s5e6ZyvfXqeg+Y8NMOqIk1k8NX25k8ErnN2gQ9m1nZDN8Rl/zb8I7NvDcjEFmbDv5Vr7qdyH
octkpfdjJoflyNjfvqX1VEgA7hh+xyCrKDRS3ibcmk22ZXJ3vxs6Ev2Q4JaWxGboVUDuA3OhaMAT
ryK8V+cZiORGY/B699NoMnyFRJzlVKlN4WZcL8UlXSkizPIKgiyc29baM6YZZJQD7pmGpLSZbZj1
tgjzd5tTmiwWS92F6VuZxWec4HDnZ2rt12E1C2S2AU1q5+2ZUfgoeeNyqrWkhfEPD5ntPKWPi745
0NZ6d7oYU+NFdy2/vZMjkAYbxUszkwMlUHMvJweZa66vP5AXeX3cSG3RhNnRtCjS12+UkNIYUvT+
Zau4+dEM/iEBP21q4a7MgP/Kp3/gYq3MgB4ZiiWMlxgE3cTpPUJNRDoXMcIA6xkBwJ+aHwDPj3fU
Y2KYd36975GBp8+ph7hyP4IStab1SQ2VZ6iTeb4ohgtKEpAhyn9Er4z1dpPUEvmQRCFXP6aQ/d24
cviiVupyM83A2Gugta099QnoX5yXs7h6OTIgLv/y8wRTJELGO69JxPhJ9lfA1T4ylPQE8uyrbOEc
g10y75gi7eoJXDMmk3hhZkW1rfPZSS9f5QOeomj3LIPxJb9xaJoyC/NclC/I4j0kEpH1Vi1QUOeb
14wyn5HVTjpQj0je3RFzAxpTIVmVHH28lMVJC3xoZEsJXM2THJFYsyET4YlPY+s55+DAIz5lAu6k
NdsDNdPRz5LOgt1Gz0WodShw1o9ILqR5wOyZc4AH/4gum/nHZz/xPTeAw8YynXGyW+Wfpl/LY66/
ugR5rVGgTM9fK4bfU3cftomp59dUblw/8FR65xA5pnuDZjvOHV2wOgrpjK08t/oWoS3nUw57hVgs
h8y4NW57D+aritBl32cqtb4i2c8RLcKwHuwuzRJWpSa7fkjvEah4kH1VdXfy1iAIWvsTpjWjCR0R
uzM6pVGLZDGqbqSbv8hmjXzu32GaqYFBq0pWa7uLjyGkrRkO3RONzcCeTLKs2PelkpYg7gZJj1IP
4+1f1v4muLD6VLI/Zo4EuCTBSZ6wy9lA5gOKjCPwDOLfJslz15fCDq02b3zqRQdRTRRRkqHFD6XC
lKv7bc+fvbvz8N8si98HMXVmU5yhy4bqSrqEe5woEJBWLaO8TQO5NAkLFD9xbAP3TaDZc7kPEy35
tdRjDpsNWBMP83Ln0xJqKz9r4ue1+I7f3dnOQDEyA3d8Th0YX5PZa6Gw8qQtTEYoGIqsOIB2RTje
UVzt2i2GNv0EpYAv/vof/PMgZ8lUuuSBehfap/YTofwT8fiMKp4QuHoLllvulDXgVnVlaaw0WVRQ
xSxkW4lmHkJBg71AYy+dibQ2gHQBkSoyzJOcdi+cgVcYL23GaGaQkybbzm55mmmo7egjzG/0K7M6
Fkt2CkpiDwF+9Hd2CQX7+BraEQrcGHPpDpe97sF7Cw2ULSBVKje6BoXwRxgWsREZY+Kv1wCWirHH
IzyCZpChjQHyc6LGn9rI7V1Tg7064Pyi2giMsSrmyR6oVm7jsfQ+IZstWcoox1gK9W5BQ5b5sYgw
BdtGeC4XZ72tBVnxZXMMWVa7wbm+YUGIcl2103l7ocBs9MjwHwkedYJTamSoyXB4o++YMQp1oUf4
pZ/Sz9Ct+1Md8uMG2BiEplShFEQab/krFpuvvjM5gY9dhhB72GAztsomjjJalUDbTeC/GljS3aTO
wwFzBAcbnPvNPEVJNEdnZJeDWVRvofsWMg+I+uWqvwIujTWDXEGsJ8r1nkVK13dYGszMW1ElsyeZ
FKgOmwq+0T8p32hBqiJ5DLPTjVcUmL0E4QXcszPQoyIE/8fSgKXALY6hgWU0y/X4G6MDhmitL0lz
BEK0xvC91G6mE6R16lSgFygO1nXjMU1numRDYKwKVdyBijvy3e3kJR/Gx1fxN5ZnrwYpN7dHEbpl
xq1yFSV8wl32UyokxLe0fFMjA9EbSOrBpAALbdfYkLRQ3TRTzefCNQyB/gI1H7xVHQD8Jy7U4r1j
RfbY6Q8MhyCWXW4BCffd/rdexmRi5gya338rIwZNa2AMla4sBHfXU/I9U6oOY92ua5WuQOpq5xmz
S4Hv+Pmg4PcmvspMHTf0kcH6F92pNZG6wVSylDItySPIgDV7G02VSUmj5/ry5Y3tmwi6/VMZhncN
pPVghRpBlobHXtgbvokdJAd8Nlr4SrydJchgOKoe4VegM+WmBHS+y9eG5ZrVUIvYqFX8vUTKJNBj
0JVN564bWq9ruLF2ZoSbhbH0XJpQt94s2lEsN/LYZmMLWdJhVyFyHQGVcjzFXXlUkaG31n9a+t8S
4VcdW0cKzsRHlyMMTvqk8UiTMBbF7JrWYAQ/EoI9rLaD8s2eMe8iwfIhYs7XAitlU6cwn7+6XMZD
Ci08uf7T8Edo1UZFGuFelRh5ofYWW7EuKqc+aAezLoDlVSHtYjFuvcCzRQ7m7WCIUkwVpbtToG76
+ESzZpwCH3UcXfJEL7kMVaayFEjhzH8B0+FejYpa5mHOFncQnxVffVwkAjzOsEl2gbCpNxdXeE1A
qGV+vOQD9R9c0HBRd1paUzstk57XEayw0cgi988vW8O94KQPRUO/s4vbuaPMTjNOASXJJQ37HTiG
rGCkWagiKGcZuYF4G3o/CWloF7Zjd9F8yXJVUiv6dj9FAsjdN5D/KxqphyIOQXypRru1/AMjLsK8
n2zVcdShmZy/ydEUJ3QFChkn0/EONHCfslX6fFp4A5h+8ky289RbDA17ITkcDxfsdybUZahiEhdV
SpMqOhNZjb8MTgSXVZbr9L3fHx73A7y/iCLeOD+YyGM9GC434wBLRqNd1cwlgpZWGQbjyltxGRkm
rusXRHyioETT8MPhaqKw6GwUg4RvjP9upIVc3kcCxHsT9lcnzyQ6AiX8/5++mEYMlo/TlDRqwC1S
DTd21YstiaEuAoZ1NdQEsX2tqnXFZxt99r0KTD3kYuTLcD7rnHl4Sfd03/foSyO421gQVEja5ihY
KXQBl0e0D7TaI/7E8NwcqUdjIbp3Mqc4Fs9z01+Qk3NRcDAK/h9BSAI1Hm0636wQjEM7e2wL8gRP
TEtnmvLAdLIWfOYV+r82yn1Z4jMiltv/lfTWDaRLlQXH4HNmmy7ZdcfF58+IEuUtlquksHeIHG5l
mGMfj09HklgyKJ2ZDHEAIUlHpHkMPx4ikSLR7NV91sDknbd4TJ65W5iKrWgpkfkZeEn9h4mpc06m
mrkAam1jhFsJKQLDODYWWEewwVEeBBZreSD+cWFmj841EWi+Ha9JNr6UKZjXtxVmyEdTYzAwXce4
+voZx71S8ET7GdtQn4B1U6SYmCkJegz3Lhs9nH4o2wVJxuNO/xIxS5Drq/mmyvER+EO3mSNdtvaJ
3fW5Ql8KLgauEE9eGlKcgbEzj5K0yBDN1Y8Et2pteY8wLbeO1cZOKh/vb5FXsCBWL/iJ8cWP4noQ
8SPGXYN9Y7hlSOXzljG5gQh5sVMj6DpXby4UfLtKPpeyu6Fc5BXsYwC9gw4F4CDmpAEMf+ayCjlD
Yk8VuXtmqrIEHLf/1c2smHPPZoYQ0oBvvSS/ujAPc9EfLUJNDwuwFbOpOqWYp4aW2SXlFBdSMHY9
yes4//UtT3RD2Bfyn6KXSmPo/5Ew5UB6bD7MqLVUd1qtfp2ztHBkhMVezkYcdiGj6u1LuvFtND6J
S5JPiAPTFO7MeVgtL5aTCgc5xPSWnx8VUw7HC/aKUKsYyuxHU4ghzjhxgRw3KcGfGAnGRta/3n1U
iUMl0AfCzeehprF0hDMG9+Gyn30bVrJqga7ulFdCWgF3BLYG2Yt3XRp+ZHHSE/BHCWQUehW1Gmhk
fc7aAfh7G9WmysSeOqmfDfPlaPTG+8xBLa+GW5MXFVhfEdS2CM5rz+l1yfCn4VflKhgkgAQC9NI2
IPmq28K43cIJs65dLs6zZKE/YwQLjDYA/iCs1LKcIZwvWR50N1uQfoSxILqhvJjgEDIkzeyJxQJE
2g+2LfI8kFqhQNiBm2P1toMEy2xQ2N1YGzXZU2pOg4qC984Rvp1o81oBsmBK3qQBwKupU5Yw2rQt
WCIowbNHVKTRPszLm/AoVBjpWvI2FEQFVAbm7o8azx2l+I8q8DsF/p6kq824qsi/YK4wfH5DvH9C
7BfN6PiZWtKDltV/aAE5KTky0mJD47asIzsf4pqU4c28U7Y3JGTL0ghp/rMZsMeBm3htOU0U7Mg6
hXLIvk22d/yjtAO2GurVaM09FYGVB1mQ+VSmenTwof2M6JvZj54ZLO7WdxzYzEubeC66svP1OKAC
+p1QC0ztZ3f2O76Kk+ef+3nvGytbznirrBLCOmX+V5KYyDayOA6Lxf7Jt8HnFQdLKVoW6CbPAQDn
5Lzpue+IC97U2vDQOn5dS9BxwWfrPnQChMAS3YvLFcb72Fpc6RFPjS1PsC5hHpgUUt/TDodGAHuU
H/n61MPlDl2lUZi8JmD7QtO7A3W1v57s3J0Ocjr2ATEgTMBh+1HA0CHO6ELPX1zzCyrAPUli4L3X
fNfUx8qHwBb9DHgfLyH4vGc6ptBDY8qDdN2uextFTV+rTMzlDscHE3u+wkKjPtWJukf7DW/SWj2I
kE78r8xPcQ3pOrPx5ihbLzo0wRSrAqnjqj8h8xLq2r+jM8JQHO3QwMRkMQ2NZqAT2wYTOxndHqBK
ekdQtOESgpowZmgGIAwOpi0gA9vnpvJBuZ394PHmkQfl1oY12oigW9ZPn/X7/rRC3LJPjSDebNsL
ahUll00AXTyzxwtHdfVkHwNil53yex3M8NYaLubCqyjGoX55irejdwh8XPIDrQFibNP46Z64WFgc
L+oyBUWZD5k/QMuh5drs6CMQ7pFpxjjx2liYks41MOyEYOIPp4qkl8iSZssEt8foAUGbjJ9Wq2Ol
iqZxSLZ8rHTt7EIxWoedG8Y5doOkAUjnWI2KUwL9NArmJXka+ECB4MpbT5fx93Ht1N7+xo1isAMj
wdXsZGYt0BuowmcySv/o+fXJhPC2+UcTXJBiWJNqFl+UiY4Git/jj9hzy6bVE2AoNcj1MYTBrVO0
UugllbbGjGI4O5afGzb61yQSjyx+OTTTPgVslCpV5+DpsC0GZ0Uu2cLeMbj318R5lI1XQ3JBOb9r
yKu/1Lo13udO1UN32ybBoU/FyczCCPd/2eieQbReacz5pvGQvvOWbxFHd+tMQEZJs8bJgUVFnFNe
u588dfARK1e210fvQy0+X2UvlkADC28JjlYSHebbXVXVoVHiSAXP2FA1UhVWDMt+eb3h4Pb8MwGB
z4pfa6ipuyVpiuVnwt1itUdPj2lT7anchIFRWldmbZnp5gjpYgOrU7UplUk3MbWc0vFhUS/LbW46
YZw+GdeJ/yxPLPBWaB5eA5e9x09j4iwR4JUey+BFYF5I6HcmPf2QETO9Pgg4JT1zCVEndzSMe4SW
qe1ufJDwhFSToLydYMFCqWNvjabwF3wUuqqOG3JIk5HT7vlGzsHb6+n4pjfNfALEYDuKLYYntGJn
miSDYSpsxdTxGpl9Z8m88hXhh8cCZ7dT1Su1uOpy6qc2FzuCfe9u6k5J3e2eBXBPubG/e3pmit9I
ukPDmRnnWfpgcySAiqYpSFJBx0Vb63axBNX6Zc8/rP5OUrzYcRqTkbDIe87MQu2hvEAUr5OeP7Pr
4othQvldkRJsowPfLE+uUmLaq+9jgfNVsLHuIi8GAnYGlbMJqKAcW3b9CGmnInx3JKR0OBPSj865
kpa9vn/cstuEtwwsl6z2VfS6Rjy94dMgQUzEiobmgu8kaALj19y+GQPxEWg5XA9i1TtLt2lej+sk
pem5oLn2i+dXKJ1gEQkXM6LvZtS13hhWKHWZ56emN8mTl3TeyouIVaETDQIiQbmlB8y59ElnU36b
9TKhf0mS2TydANoe5LQY58IpS8aTIjPs75f32OR62cSrrmkXmuoGjY3JbmTx9Y9pfxqSMYxLc4Ku
IHiLpNOSfUCrd9vvgVfImOOiBIpYAU7riqT6dZzbDvfjr9TKSVDAXbutmtXIRnVaRV4k+8HGmdCF
30ChnDz0JLp8+IAfmhgV/0tPhhgBxK/yAxNyKRGe7OIZMawwJsXq4dQnHqWKR/Etx/5oTryIA9NR
QucJ3adoCYwbvGcUQ1sAQsF2DcHGh9iUwVUjkfirCADNWzEmoyExUW93wNPc7yV0Wx5pTdGBVLNP
C9TAT9ukaZRpJ+HowxcSXRycyjS5VdR2NfW6CTgvOy+rszDN56Yg7dM29N/ELCKIEU/lMXXWFb86
09SwPB2tzyMrE5oC4iAkQ3hICzvXjdRUJ8xzqTwejrPpQz+IU8eOJnKAeGlqeEhOssR98lMryLSY
oRUHGkYog7QtlX5Nre3+OvmJ20+5lQ4C8dtefgx+4z7KhlbQOObL8AbDSlKDnmNFVnD0BXabwi0H
7xJKKmSIiqUfo2X5waIYyh8SyCNyxBDXKV6T2c6MMYXwnCjXyU6jDYoJrQBKyimt7HSpUuCVAeRP
akShd+cN2eXBQxl1rELnNowc3x093PLJqsPSKBm1n8ehd7UW0iJwuujr97AX2XyS7PZjuUp6+G65
zftJ5mim4EE0VDvqnkAiK4+UXzlDrUZ/L2RVeQpZW1iOWKhcLNmFw8nxivcgTei85wYdMkKqN1vx
qXDDR3wydWwrcovmzpleZ5p1LxycNjrm8g3Fpm0s3tYaZioChMyzvXLSMZn5Z7mfKPRokysodz7Z
TB/44Pn9hSCR5TewDC3yfDLnkcG1BE79SES8Bz9Q3455tIy2jHYJc/l/0QaXdlG1gx7fnrNn55wD
t6c8EMsXah2eCauxsOAbf34aU0La/pot1NXBMLDvFm6igFqDLNmuTU4+ZE1I477GwXwLahJKbX4i
YypZrp00uc2G1cqKvHuKy95uYq89RBTM2jBFmFZkb9BkKW8IYIC72E3c03mvXbuCGMTC39UiqnEG
D9R6vl3yQPDvWxXhkmCALuH9y5BRyHoCh6Uq8Q7lWpWQaw8AN9riIhcFBKRO1m7L55jyNLeXHM1C
zOegbmmsbFachKtTkRKNeE43ms25t/OgfNIJ2A3SNFn5keineK/fYXeqlZ7z7IdSQZHkf4drlLQY
OXX0Ra2crHPINKtGJEWmZAGvjC+d/WuYiFcAQ0bYqHNhMNZyZnihs/1O99Z+Ijx7z9F9wW5hvbFD
pfkae7v9jEu+SEdkBZ9iWymhJjPVrYk0PWmCCs75tiTqr8cumd+PcXrDjlvVtyv+sq3g6Ro+Ld3I
1w3zy0PUSEHQyPzirH6zo5PnxDVQUtfc3RDVsDgX5O28KNqKMB/lzrjIrnGaMjsayaTk/KxNDq+p
tr/zRoTQ5vld9cljjOTfzNiN+8Vvgam98W+x46XVY9JWVouAZsSutdQM7ImLUZc3eewLaqrPXlBk
lfPgGQd1BCP7BggsepY5X4GftnQpsMzJz9nl20Vnrii/GVp1IU/HbOGLGY1nKThcavVII4QbV4KE
ZL27MQgICAUPhaQPPUlymOXZNaqbYQ9iXh2BA/z0uLwFbzRxfq7TZefpvstNkO0M8f/I5EABAgMB
NgPiBC9raw2sFd+wZCi5rWl/HU4rebN+Jc48qJoRq8SB/nMBkjiVmljntMefvNZqyiKfPkSNnXDG
Cx/iXWoL0r6uz4L+DAOeBURjG3PnNMzHcWe3yy2cFrrWpt+lQhLcDdnYfrxBUcATo12MkjejPCAt
FpZdwenbobP2b1tljqeS7PvP5qweLYBGKI7SkN8oQrCe3mzLmIW3riU4IIqc3bcaT3WVm/tY+yco
2Yaa84+bb+Gh2cjvajQ0g44Zj+rI2dxJ6pmvg8TnB8u7+quCj+f0oyQRORMh62xejAdq6x/WytaI
+5XRAZ6MlLA7jZ2nnFQCr1LYUEh8gJqLvvnP4KymeydQgNpwFd/qEiawVcVfwWTQfAqOHaiv7t0w
tGfUE1QDZnkIZw8olRvp23lNh3bDwBxTUqcmneWPbLYuCT+ctXQ4YsqwXNb7+E636nipXLHXGkW7
+ezUkiMKGRyrioUNkuNVW9AcW4FOsECKbsU25K4I6UQnmHHjkJxskgCt9F9md6/eA5hdJhYLVRaU
hFpPPRvc5aglwxS+iwgEv/uXUx0r9EFSTYwrNa5auSlv3mFtZR0lnvUOZDeD0Bpk2jkfn13wtgWr
T8PXYrk1OidDcdA+SwQxHxwHfmNnNcVCOMyQYLDlEbY3Wru2/MLb+8tha8gv4LdRTptEYT2Dzo84
IlsQMTYbBGJ8RsZitCjb9rRvVuH596jDUfSs3Nplg6H6aGI39ovs8eeZLosJHnKbsgwaJYEhDnzC
OcmeLKaiu0RPHSr+IBtOvvQSyHnaB7ododiUwu6jcdk/GQvNyETiBClOs41FFkVfPRB06C57ksxx
q+J9zYSqQ2dpWfOLLowF2mX20HY9SMFfnWbVl24leIhpEGR5pUqOSJ6w5AlRWlDhiVtsSAjek+zb
H8vN/FIgWIBdCfLnBKvFSjZeGrdDi1u3lTcZJt8L/aBzjMLqmF+EqZOw3bxGLQzLQdhiDxtHmxxh
E5C2MLKRj8FEcr7PPD66UokB4SHS/qQhkXujlOS91D8oF5eKeFMuT9nk5p0+2sykkXpTHOS/ia2L
Ltf19FcyCuGraS28jKyVZrXzUYDh5Cqze09Yha1KIj0J6PrI45eQnqFmfSRvgkTAMzlpOv55ZOQ9
njogD6mG6AqhASAAJYCbSyUpm3oEIlv6e2kbpLTrU58fLOk2jngYX4AEsQp8rlzSGdLEUvKagERn
BGNBm59KSUKTeeWBDb1imPX/X3Tv54cAzuf7Ll0ldQDDaj3s1QJ2JBnjrj4eyx8ExgFiBOQ1JhSY
0hVEB0JVjA0Pwx9dcLPtQy/5tlagNNb85jkU8dqUwoQ8VwPhGzfYS+kSgH4BtkDXe2SOxMhLoli7
veZWBYBvaVOiD2mdJ4i56mgQIVxnMxBhSkKyBMJTqR73nZrmqI3WNCBILK3TMQc7o/IcGavwb/sD
Cdgw7fp8WsR6CndiZwtTT5BWTl9RrzHlOIQ1oXeGWXpFVSaMF/vZuJ1+cykWKjqhpRwU/Ib50Z7G
qMHU93v7qM5Mj65lW2BJXAuzBNn868BRWhf7Nxwpr+qCPN0yn4DHAJAbaca46JzF/l1AUTrh+6wC
61k0WaSVf046XEYvbdqzC8Mmc54fuIWyi3yn78CL+b238u/W1d297Alw1xkCJCTjH0Qv+j0I2Zh8
KD9xfHzm+s9WRyK1RvBu2mKSwQrgOCQLd1nSiGFvJsA84ayGOSv7RQViW/oaJqItzQg+vlHaJsdH
KYULvL9NcjYdKdcQkwFqXSXSLyAD69dsdY7IdRHYOwtmgApI3qamOFCjaARUqGblquw6UM6yW4Yx
EkxNLgucMXyLUsHNx9OSGDD2mAfsBE2nmLnO9AkX6DOCkxnmNUZAU5q6gBffIBrocHXqZ8uP4j06
4XRs6L6u/uTipaRJtdT8vGys0A/JSyVXGWI+13fjwYQAPrmKA4/Cd+13f4pvpNc0Fkp1gHX1v+RJ
zMbD1K16rRlK2tiTjHlZm3NhpPaKGrBd3CNepBrQWQ7sRF+WvJUyOsFfgzHUA1e9uoQFOYcz2gOg
RP8M7tFfLINxIE6OAh9QstFMfocGZk/T+tlKQdmAQWqW+TUCTboHhcx4yUWXNshZyssItS3rA5Ib
J9BBp+hNcYkehci5My+PT0j0ULsTH8rrsupO/qK81FhKW4KHLH1ygT2iLR3sg0urg2U1CvN3eveg
ahnfGATYCO7tu5YWEOa+QoMfZqwZr40fFAyodykU5sphG/9zPR15CiJQQTaAgf8xt1e9xfqwhwEz
QbQrEUy1553YEkd7MNH0NCH/6xrGJcveTvL9jZu0LojuGKEajVvaowNCV1UeoXfSU1Uqkxh1QmJj
YeK2YKQcZcVOEXH2UPBYytoL/H2K6fMVoWMTD+0y+3QvFuT0qWgRP96E3pUkHA5tIG4VXirkWjSC
LOZvAI94eNKdGx3vvdB7dofckJiWUajFYxuzU70tTLhp8kEdiNV46M9nzvlwJjiF2dEIHhgJnl/O
Viy4oB50bVaxVICqMyCAPahdOEAZ/EJvbJJzeoB4Jl/025M8/JTzzqZ5WL9GSUxqEnLRSzfgyON/
ehyzI5cxTMGWbuNX+hCsBLUA4llUA9VHhqblL4HsqQh5EULGENYMrXP9HJWPOrE+MNLbpMqPvzMU
BazZjILg0t6fyAtgsjzD0TFJEdL66P7fwCk1D7L4pAR/eGdaNcvETM9n8Sj200Xv0XxtcMburK32
qdg7Gxbxw0zozdF0l34IyYtqQSM99oMa+C4xlHbQ7iq0CzCmfjrD+PXRy9ekKCpp/y54CnYnuH9O
idtqdBlCcxgvjqcqQt9vhC1jXPmN3SexEXq8qd70fvo2rHrbs1ZTc/3t3NOODhCMwKEy29HWQ/Pu
p06pzCTz0309S+u4fBajLyVJRnrqL5b58SnkakHLR8zdAt1Kpc4DDdTVbl0bk7dwhdpRBdJeQ+HK
rzI+SPqFvWXCaWm3/fCkdgzAGlWHXQk2OfE925bm6BiRI5luksjjO6TVZ8ftzJQMlHMsfDfJg9Eg
cMGAHJp/5zIHH2Pb0AzNFirPt0dS+FXplag4Bp1wCnn1bGo+sMjzuLqqvrVp8dmBcX4CSRQDB+7Y
tY2InnoSaugb9otAuHSLI3wuiz3R6cqpIP6vfVMDHGDJYOZhN7nS3HrXRnQE7cM6orsAglVEC/4c
Axi3TNYzSU2NJoyHd5kZT50m69jYX1wUoUZU+h2b30paFYujDbSqhyxeMTcJIWQaaA4bZ0uHsWCG
R482TAeXkYVfhNC7WNvmcO/cALIb/1xIOe67tPk3+EKysTcCJiP1u0sKkMHaOpV2iDDm7XJWL7MX
3B1LsWH4zuFHozhY6O0twua1MLsoR8KYP8VjviB4B21BPYVZOWv9DehfBGsV+d8T07b2q1IUSPZD
Dr8+ES0dPyPlYV+L81FNRZjnlxK1eqGDL9x2E4bbx47vJsa+sjBLXOJCcEhS8TpHqNxQnmmmbfn+
tr5C3vLbPumTW4dnocm1Rmw8IGtgR8PzZtpiimfoBoyM8I0VW5Oa8eGeFEQeCFgIWKE8HwgOEHkY
W3C7Aj0SYVSdHhfWSsAI2RQ2k9hodZYSbUUaIL1vsEocuMPVRY7TrbRyIBMpFSwl0e3IYQ2eqk+F
Nj1/ytkrxnpx85rZ8p+ELgpfMvhf7jUB9vUYTfng9ikA7GU0P/EfrZWRO7ZHW1AKLT7jSGHSLZPk
o4GUkSzvEVF7qPmttaPEgiHYDAK26ogOO8+NyCJeqvv+6+MYlPbY8aLt73VC/Iog1kCe1Mz+I/Gm
GMs3R2oY5uTuZx7yqVhOSiFQI+NKJPMh26tjUagpwLjtYW00tOLfGWEoOvKey+8lJWKUdiaS0EZw
DV6kvCDDhCRDcm1tADDbo/sz0KR1OMdpBq2HGxWpM3fQk22plgM7HfcBwGHnhv4O/ZvvRd7CEhis
vCgy+iSHQ5z9Ny9TaawCugfh2U7gmF37JuRGLcQMqISf15DuNRPx/eDMPnmf9FxLfwVsgdD0YNYm
KY2nQnvkPqipKRPEpqJK+X15zDesu7uv2NbqihA+SE1+wQ0r804NXbLp8GZu+l2S4XjqSkBHoe6Z
I/fy0V/LGuXm6PQIZnO4NZDh3hBmt2Em7R5IPEu1T1Hc4mweBsI/iHgfjVGalFQ0ugpXHAGGGPDl
GdCebHyqCqDr2ZsgmNGo/GTeYAeWVty/6estG9v367kW70UMFzDbrHQjThpeZhqxNYYQU22GQ/Ka
Xuo8N40yC6tl2auWLgr6zFFqhbB44Gba0WVGzbYQpExCLq2BC26N7OxRScR2IJNkja4HLpTHAkZr
tSOWHlqQbjGvl/iKCHoWqrC3u9hHCuDkFWeTx/EG8SAJUZ9PW0j/y+0bqcVb1xI+q70bRdTlV9IR
ZpTuuC4dNvnlw7JJ9Qr0HvzJsCJiW/MaOFBzF6+1BNH2I5iQsd7ravV2ZzpLTVPZui/il+pXx3DF
+7yEYw9af3/LYuZLGwUBR+PPjqKN/Bu//9FDHQoXvejvaPNblX2CJMSmvcD/JY1H66UlhVcj6VwF
yqBENHX6bj7pgQ093FL8OVZ/1s3Da1hAKoP0CY7ZIEGSwCveDO64xqjXSiEhEqcwYCKBqDSIu4Va
y6uC3KirPDKRXyk6tiNWz3/+voQMt6/KF+nuOhwr0hTYDPh+F4OTMVHywmU+Fnn3PIItCvPCIPSq
dDDF61hKEJVINPjJUgyllwTuonc78xFMVHbk09+76oL6h9QPKI05c2+yeX8v7pX/0ekAoyx38LCY
RHrTpxmWhIBFBm+ISZ9U8vVzI+wq7TqkDablPPWDcVcheWNT1wBJjv9+iZMlrZggIaX4gXrw0TRp
GWWr77CBtFaZMbBXSoqTfTVcCx/VWStgyV/YzBe4amPh89YsUA4Qf/h+gCXPJ5pcBd0zh2YksMqC
+Tq7QxDO/5+HkQTjd+tL74Pi6n85AemYL7F00Ip6ZCREkXulLj0BAuRMMVEGnjS5cuGYTniy3dlX
o64qKuYWM+kKzTsdsJ63E+OyN6TthytxeNQEd3K3kMKRGN8CSj3u9Cg7lEvERa0Yn+3NP94m3AAx
aj2zrUzidJATu5aQyNXtNpoYDVBUo5Tz+22eUF6xrngs/ppjcLuqN4z1uiBL8+Vt+ABOWov3dRi3
DreFov/qhnYbYVA67MsIcLE5LK06+q9Tw8Ig0XKNtLTsKXtzCthOrEi3LmUwZvLEmE/pQjwvEP6l
IY3nyRNg7UhB5Q4ckfNOOtP17A2HEcYk6F0DHPXJ5MdBrw0vTxjFjDBT2khk1FWc3/3YHR71VorL
Y0QFweFCgR2mLpgBiEa9Slwu66v+WDs7ZlQgrKXijyBTz02ynv09ac21GCY3zvySaOisSiqjEYI8
nlqvJnSm4MRVbo1w5H2dX6O9f2tK3bWB+XOxUfjMtUSMtE+E+8QBOoRt3VbdR5qyFI0tXc5mbX/6
lTDiMhWq+Hpudlz2RYlOUv4DCrdvJz6jNCJemTuy5agquN9jLCAEI3QWhEGjBIPfiZ2cgDokKbGv
tv5UWSjiFfDJHTh9NSEZwP36Gh0qlBKUDxD8NbOueqZecsi0E+oNaPf0ENi16W3UvOBWn3cVfhuf
XeKGWnZpNNuwIvuwlypSpEDaw6MiD/csTuLYoUJs95he2MlI71aXIhg5VAqV7Rspz70qGV5t4b1a
qWkdvwEQsw7xymKq0dbtYwybnWQPn39zgpEDkrVRlencyVJLwQuPbSj1dYlNClv2vHYC2bhWNha3
Eq3ftyqtbsSTXTDpImnQp3bunL0y95QdgtqqwM1DKpzEpd3k0W1nF/jvUYOhp4mIGc+meGZ0zZib
ffx+tQLa7Ihvfi1sfnQB82cEPIQUr6vDvhDN1BqsgJO/yOgUkqzDt18N6diPh1SLWVj9dzPKHy6y
Pc7dMqkBko6DDL8RDovMag2XnpaMGeZpjyeFxi0CxL8JFmOUzU7Z2qDSJ3EYnPWYhDdSjEDq6oLk
Y2J290wh71NHpBQpaEfyYCQxzsgTYHJ+5aVgJdclnlcEd2p/dCeWFCcb4E5cZf6zdv82THAZu5vj
Q/EbvORQcGFaAJsGvUz/B+/uqbGkhY9YplSiHRAWmzrweDKrqlO7NVHJOUF6d4kgvYuzmWuqmaWJ
3BEG+TUIh/dqokmYEpJo7MAXChJwK5u7+G/0R47WVoJ5WGJ3rewO0cIqRRDSfAqwI56kLweOJwuh
7yD7IOyrcoxH1eIfHGOPktiRTOc7L5/TBMCzYuK8wyKG62BEEtvxy1MkJZJY6tjEsb1i/J2EGFXT
6eOMktDJLO6vACpkgkqTa5S5AoxX7EXSm0DQD6L9TDjtwE3pA2rvc54X5EC7o75Knx8l9fOQfU2X
FhHeNr9yzqXiw3HS+pWzSaSl+T6aGC3GVt6mM7l3tHX01xox5ioPhPXoYXzcvmxei/dzYEM0XqQN
bKkGl459JUtlsflUHloD/OTI+u2c+DzGNZK1U0rzBbDqg8lmjfS/W847THmmz832oRo+7SqPBGgO
8GlOQPWTyWnwuq0mR/a3Lz3fv88EY8pyxL6AcVkSGWvPxtGCjq9NcgzqKFNprsYHm9niotwgfOb2
e2g2xb/8h+nN2hACqzghwAZgG81lyJmydfPy9lUZ1cHe80iXWGUWDzHYRneprotTJH2bjcdGnOQ3
PFldN1739RmLf7PVrA27xqy7raYSIXvutoWfcTPTdxcp2qoEFptOab/OFwKG4liFsyybg/pBtYAl
fZt4+U7y274Ibl8DR7BjAg5FkF8LeRUujZONzNaVeQnNxzFTLzm3vSWhTMKi1IsYDBtwh64JCfSI
xLoG0o63omJY+h0xRqcxfQt551c4nzSioczhDDmlX4fjuRmGkCQ9lSgE4IEZKuyf7O+Dtlm3ESoI
FmlmJIGqhj03Iu9+wxaqWE/JorrAo+XN7bgbfrKaK5EMyKqWrTDMv7+NAtxeNXjTAlIdgZ0ris7P
lbA02iOfGlC6RTmQbToQR5sf9Jyt34je5yZp/K3JYeKRTvmBdhKlrzn1CJWLXcbsZZuYKhxEpwb0
xdmKccceYyWumeSJA7x0ZtPLU0GcyFg+Jj69gD6GuPGzLBGBsqm4JuMsTxWkHV5Q4o23XSyqO6W0
aP8IMRTZitj2C87QPsI47ljmrlLib0cD0BBupmaZXfiAhfSAiND3kay388Ya77D8LQjIK4VRVjVL
yNhNSyRTkc2bhG0/gNi/4t+Mtr0WDQ6KVuJ15jk1orWhcXqyCDFpe0p4IxuWdLWn2We25SIu7JzM
Y7PC8UkhzMqbeLwQGTjBmq7nHOcP5FHUfLQsA8GEf38ik69ynLHFEoazLpjuVwrHxg9cV9p2vNx0
ogz5SH/JazNq6H+mZ4jNSolEnMKK6TwXgjej4mlzGc62cxLV43aXSmfFKH67ZUj/somYSrKYx1ai
SKBnMOh5IMJ2/8/o+im0vfk0cy0Y6F+B3SQPbIKW4fG9aFtdwBzFw88rhT32BUa3BoSxquLVPkxJ
nQiD9tR/7flls2Ru4pn9K6f8nxAdi9tI+GOBB3LIQIO6bHw1hnYg494NjUigm0ICgskh98quBA8S
U43vyZ+4hiZRrI6NPngPAsOEpbF5DWobbdNdRUdQBmkMqgVlP8zAeZSz7jae1+FoczRpSnSPiyz9
cmNxq5QUTZqMFGlJreGEC4uEkAzBsL1Y+XAK4kcXaAJxuhWlBxf0G7s9CJev4SWU2BOegRyHGkdu
3QAc/Lln0NfWg1LFzE/8AxV9NYMfDw9TPMTKktWV9BxINXQOksbrkAyqma50c6uDYrqE+excGjUZ
xiy58HXSU5WwUAIXBZPoD/VRNLdtA23KBb0HB0WbrUvpldagoBrF3oiGxq/5omWmA6gtVepfer+l
BMH3GXN+ijBCpHyem7WpEEbAjladme5heZazTeJn2G597LTn/jZnYL1jo1U4oDFFcIv6gR1hxWju
ddGwhJwS/2KJ0HC/wItrQdR/vyMDYpTNLCGSXRCgd53NUF7HhFfw/hGMi7Zm+bsB+sjNxdYT1nFy
WNVG5icq37vXZo/3D2FKyX2qpIueJMcqMeYvkp/MXBaOXenW+4HOzVObOSJnza25FCpkSWZMAGJn
W7tRmc0cpKT8QnoPRSLsrkV4ipLo/5mEdguqdFDe4jKdRf0Tl0whjZjfVBAf2TMjUZCnjGvNotac
RkfCLPo6W9YgFhFwIcfqMwJel49EcOdWsUe4yHF542fxLZNQLoe17NWZ9GepLsUGTlZeC5BwEuAQ
W5Kuu4Qyd+nAVgacGOyZQnrW3y4cO52aQ1WmwBKcyw6jXlt5L5T9yWum/cCuaw/QwgXtlOteNx0W
yn+SreJP6r24AV5F2CzIk9FEyxbdkp9iqkuW2L+JVWGD3ScWnPZI6frSShOx9T8ifKU6g06KOgQ2
DPoQuZjUc4kbjTpD9BUXRNlhPULOUxwo8t111gfgwN5ZsKqqxqL5WO3y5VeiP6LUFWUGFsdNHU+7
eRl1A2dZvZPMnKRADMNBYSTod/zkbXxYAZU0Q4g3RYL8NMKWCrfoAOtGPrRY6dewmRc1buBNay1P
cW0mQCnVs1PDn5cYCiN5XYajJ7EOHc4SY7ZvXl/rgNKCU7PzRqOJNh/P0Jz0o7pR8vWL4x53vq0y
F4nco4AMiu+N194aaSP/SALTDGV4ku9fV5tN+X5wx5WG6bzC4KpxcPYLZ5f90rl+lpkVlujklUad
myKfMdkdt5T5XlobQ6oyy4nA3/WyhNodJs+DCSZpda92K+f3pzoUlD67U71eKFGXU1nN+sIkdkRi
hdwO09OSscWT6XpVTk0zY9Nzh49PD3YMxlvOWZC7Wy6OU4TFfTwVxQfXsrNwlb1r9AeF4mBq9gzi
7WcvGpQnP/DdqrkKOKqmUCvjpqK+/7kXaMmUZcV4ey+HPV4T+i2a0cMFB/oP1iSWWptN8Fefi5dr
R55a58YDeVkMsgRLMxpmwq+OsnRXPd7i67i2wvXl0gFv//nJVMDCjjSmis0ePj+2d61aGXxe3b6k
cow+wByRlL7tk740RNB7AV0M7JVeC09d0BI6wOYwPEEiCrd+r/FZsFx0nTX0stINOp4MixKoVUDm
x84iPp7a1LN1uI2MAy/HrHcPku4JglJojFSMRCAcDVu9WL+8JgSWTznw6vxxWh574t7sILsv2d0r
LmU9trIGqjmfZkCOl+jEW/KzzF3K4d39/hKend+MpgZcLZqBkV9YbvFF2sCO5wzLCCmaJ9YhzorP
dcae8t4Y06pJsgyk3R2vO3yryCvqaLlne4plZbzXt3vPdicVteAwc0hEhDABOmlwN52rNfaNI2/g
wiJ7sIU4FkZ2coHp8NYm2BG52Q1bEwnKMSvxlHfi0wSReJrhzuHVGxUbmtSfkyX3QuHEPbX8AZ8K
vAYIAMtyG8HtdJDuwOW5sSy0BdIDVxtq1Oqi19IomnVBRXH4OYaQhnJ1KB1cqlhN3+ymzlpjYxOd
eNraUIsTsQW4o8o0Y3R0/iF0cEKpscQ04hWcjCRkFLmVboof1H5lx1zmd8oIP8MT/wKZPM914qvl
UoC4bHpHiA/Ts4XH/6Ka7zGfojIZPDZmY2kwTrap3h93O4EN/umFREfVvmINTnw+iqy6xZvJRV3Z
SrtAqJ88v7lpzmozXMbYYEXu2K7kgEE1Vk3+83MsKr5btnGSxJynFLVBfno6PeiRSadjUJPLejUr
e78NdIIDw6E/Og0Ar7jzekP047X7ai8/clXcCdOe59hZUzesGPWz9j0C5jOzwNnfRcRZ/taSKdQB
OqGIN6K530sx79Hck3wedzSDCz89bsErW/AHdN3Kx8nXEfWnIhd3rieVZF9iNgp5VXfjLW77ilc2
Gaae794c+M7gjXQsdk7hv2rX4pI8kGj4GGpXs1Ngf65nnWcGevYtKIqP1M5oWKgr8yuq4pvR0csP
eP+B6AOTJ2EJqLlCg17NzCYNUy43l0uxxBi0jf36ZJgxsSd2aLQl/cYiDpmtgLr+GI+YoGQPrGgZ
X/1eesQPfRUjBGB06nnHoMUYeg2nfmVsiozNyNEFeE8uHvjNc50D9MIH0vpsYu4NwlQzOsbqoWlG
nxtb5bHD7UoKGvfrNHn1sEkWPJ/oUzRjkUsIsfIJ3mUw8b+8CZutwbjbqG1JpEu5rRE0svbmKY0U
8Xmt5Q/uI359vC91S3b9qj1fbpGdmUavrRzbzXufDhae2hq6+u4m2dAk5ZioCv5yeO/kCqqCegfC
jraNPAN40LSAVlk2MFCeybChKVpyufb0sFQpGXQpwsD955VNb/rEHJV6eb59dYyYlAcp0hRQqsIV
IzbiXJcXg9T1nFO+b11boGKn6JOG23GuKhg2n2Y1aFOrZ9O/tYZPk9KnlboJDsCz1KR0rHQKBx9y
WvsS/28hfRwW8PEBBGbkSLTo1t2N15aeCHRObnmpdvFLSR1C3w96zNfEpCwJyHQeTta/AliloeXs
KefKTv+mtNixqoCEay9C1M6Rx59KlCxx4++DPiND9bUCo6irSSwbWeknw1TxxPNbFqvU3BBNKdsC
iDr3lhVDCql4c2sWyHBdkyJH+ByJ9HWuuJ32tDrjzCjolsScb/f2sHeSeS4P9bkgM/gJyIY0JxL4
wMUdFlnkWJYaq9nlEdUuSUsm5hZPDNjC6lehUB/+08g8o2e5iBqS3kSH6GfKfrByQ+9NTxn47h5R
By7b8xKE40VaMWJQO+gNaaAmrUn/U15nw7UPM/wYYHnrpADFEGXIQjiW7fZInG+reNcUiEKqDtYB
7VdsWzxmFdY3h02eoiy+Ox3AS2iwzM25SPLzQXC+I3vmk/V6Bo9RrCcxl3HuPxUSFjSxjcCNgzLH
2QfubOVRQynRAx72ZQfaOddVWzUwx4d4QWYjvB77HsaOPVqn30IKOXvNoxtybbWX5D0+UX9rbNFE
l4EPysiB3sTiAYYsDM3ti8ZvPCmB9DAiwOkDZzbCDeVZ++/IMQU27VrYddNqNubYo6i2Or1lBQ7a
JYcL04GxnNBpJSLcRcjWgVtHev4GZ8pWgtR1fcMxUvM+rA3i3bzkUcwFVCaw9u0kX8nO6JsuBAYZ
1lHaB7BXAU98S8o4HH8Fgb1NyKewFUCEepKcoPjcWOHo2ODHoXbOi78zcCQ/JUxXHr8xQ4kAxi1i
tQlfmns1wuvJLC8v1e7ZQmheJ8sloMUbkFpz0GRy0N0HLEEmcxHrFowV2J7/Q2W2wM8SU0FtcgUw
m9Ck+9IxC3kqpiUFXYhmAVhtKg/jyFJH5oMj/HdVnxuWulCb5SR8VFskO9IYyET++yQJnoe+ujtP
x+sjQOn3jinqz2pDh4eVn0NtmJtc45ycIwaSoZsw3RAQr76FantM29JaVPDlAGVP8HIptybT4jpR
IeYtmwu0TzxqEHTKtHyKgdaSIl2s12QReS9mGNG02yA0Lgpo+OYTdv7KI6K6WoFjj8OicXqL64OD
E59+hhu3Qo9UwdHhGsh6YyAmnanYNM0vCcIxvbJ2EAD/JWANLrUfyzstmlOv53eNSMEUrBSqjZOl
4nblwuXgGQVFYCV5n7SHMl8WjrSj9kXxVQVlv+jizi14DdrjOVMlRflk3vAOTxdKYZDVsU/U0iNs
kpCyyx6cKyGIsubQ+9b697w1Pr4XMLVjhLBjjad8A2Bfd/5CbeFab3V+8h5gIt9JEoS/5WwGzYMJ
YJBaHgm9TpXpi+d1ihQLnqKfV5U9gby7leqdyplxQDdK/ZosIalB1WvKli/dp8PGxjfecbwywERh
MLBHAQrJ2ArUHW5FByXJpXVepT2x8yz71Xnc1xoCwCLHUpXig54XDRyBjj54cy2FZZJGfLIhB2YZ
nJ1PIE8xEqaYon6T8e8U7FA/th+bw0sLY+OKft8LD1qShMK5s3cTvYNinWdoTbNl/hToVCvxVEtk
nhLTQG9f0gdygDJ1YejgSqtkv3bG7O5P7gp0xFIuToXnT2lMeq97PcENL947mydsfbbOkxmYzasb
9SHqptvDOISK0mrIt1SB2dTcV5sgLBCFYv3dvdcpcXhLAmog2W1tyEEqyfDUgHASn6G3lh2ULr01
jqd6pKSpL1vY7y8H/iQn5vMJu5JO59Rs1ZAcIskTojFKrBIJZ/57YUNmwAkPn4dyWq1av9VMyJl8
PKd0TFTUULc7adpwkCwtLqPzYsfqxRji163obkpSbQvlzTw2a+AJnZW/L8grYGZJo+r9Z7pwtso3
DSXzPnckud5Ez1PMgh5WyAbpv/U3SwZzQGZWbLKAS68Q77o1QWm1MR4RhJVI0LR7aiCunxl6vnGC
TkiuLS4wo8oSOXe00TZtBwkGQ2QMwIvSleR1ezrsC/LTMnz/mxsT9q9A7oj1a43TPohoHmN1COrM
DzC0E26srPbYEvWv3O1q8M1tvQFGRMlHbGQloploOQouXcm7TYo4i40DR3UyLM3TDudFr05TeDt9
quKQ8nLPx/CPBCddrB8Q+iSZuhkyzpYy3t02yx4FfThaiIEWODRnBzT2m112gQE3QgSI4pA6mz5s
jbaLjC8Gq1w8FUw6g+4AKBHJDlP8OFysD5L36qv+cnsB0Gu7SHLH9aAjYzn00oeSEmlzN9UXEZyW
WpHeCgxI+ZArw32yZ9axADdiwY2W1ZQhbJsp5yp1B3xQF0zTNNPofXm925ygGt/8NQzugZuaAYJh
Dcc3hj/lPx/LlrdAZKPnzxl04LZ4MBOUvDQcDipil65Qv0h8OPlJjnvMA69CBFHhG3u+r5aCnfT7
urdpjM1SuBMh3B2eX3gd06Yg0+IROc0lvZlpLq2n105MrJEvNLR3WKjceDPwlvvpHLqSj2Tbfyj+
7qHIHJD3nqEjATHdl+8U4PhDCFchR5wo3L46AUIJER5nsBtriaYnlxbTTWtVEb6k9fbJEIgiDIfU
Uo9swWfKWguY3asQdUjnx9WM5NqJhRdjvqMDmN8Q+ssOx1+3CFchSCTy38DxfcF809DmZg756WxV
iNRTUdN+sUzo+gZEpZj7V09Nn3/i+fbTahAD1wW8jftVFfnFSPET8bvHXgR/EJo6HlH8PmHaK4fc
znTqlwyUf0VeZzmYrxSvPNlE0HjqNGri42PVInm6JuKzVa5xvmZMHtvx1NaRwf/KDm0VC8qsnwLf
4dvoV/aXnk+tSMbgc9vK+kV6zBX0u4oI4lhOLl3ujO1HtdhIIFkUJK3qGLec3AHAG2vSbfR2uaQh
dxnwPbOOc/R9N3tCWI6Q1U84YtmZbBasBfi3bi8BcVdhnighazL7FtGS9MxxwsTSUpUrEnXkU/4Y
ZMXYQjadnpImn2ZJuWLeGNSPBN1qfPPkU7KovzXHr7i89JLHsdMCvyTrH6/lOOB56dFoBtC/5UjH
zGoGGOdykT+q5MOUtnpzsHXYr8UcpvjTTrD1C0C92j8YNa4aG79mrdUvoa/NYfk6Uax7JupBmxId
fGUeaC+wnzN2KlJIMdjR/fe70wrKHNZQiRn2c73edH+RFUI6fenJCHDC3CxZaPvUrBgrqz+VVt8Y
ZMiO0dwYKcsLf82d1T4RG/Hcn4rYKhAf0axyW13prXTxgYQVOgo6IoQ2NrjrMCw1JkKgky4Z9bye
5u+KgoFafBOMfN0rQZygWHcFPQLjU3wzyv6GTGkuPgnY/39WGZi4Zd2EjU+rDqYU0V7xvv6VxI7r
stkVjkVC+XZrUNVWRwycCBdFEZdsNFo7inIVTNDDk1XC7C0fy7tDyvjGBjSAkzaaypHqsLyw40Lj
TD/cyMgYYwqVxwDjym6C9sFUmm0iVuiRyn3JkAeYK915s0HocyKrI3QmUSzgtg2H4aujfbbFgEyO
l48edxw6MuQW4K8N/eB6uGYZ50O+jelkqLl0SGnX4xQYqIejTlC7ZFcbT3dYa/LNkY2qwoRPUohT
ip5zWKguSTSaH2Rz/1Cin2ov2QqbPEFLwC6gxT5NvDNlaqOZKPuHGtiZVG3OedkR65CDSkqvLyn6
9YNZzKK/MDHTo+yVYT2B/a0CNcyRGnlmzo/YkNqZsDmVpxFqMQtYuxO8Q4R9Duo0WG13tgn4qfT4
DS+hcqN4LM2JGLi/cGW6lTVY5IjfvyUDsBzk9nAmZ5yNDJwcU7r8TcLHn4zpOIkLJNw4QI1g7Ndf
RyXfAg9ZKTLag1or+pNaK5uomruM7WyWZ9FpvoD2OiQqGe2B5xq4FF2Y0nsaYMmBKeW+iYdfVC7U
815Gp001DcEFAfUz9RztEfMLWJN0JOkShJSSKur3ggYFCpQ5jKMgOHawMoxUoIl3fb9VohdQxpOk
Z+OTRd8w5Jz+cx/ra8TFQubmLsCe1GxhaGOKZRAGIrS2HXRhRy4N7z3ocRVmDG8qRbJa7LI+QHFg
kbsJtpKZ4LGDHeuz8LdQJiZexaoV2bJqXGmjJIeJvx2ttTyuUCQZ6L3Sza+0cFNCoqw5Ak5Ui3iz
HK6X62FzTGdzeZ4YKa1q1N9s6Cw6Y2hB4m/evSD+y5fkNFDw/Oqarn/+5opYcouZvOUtit/e5j6N
5ckkU+3t6zJbZXcVdQ5ClatOt5/YRkV3sm0DMSI5m1GiKDprA0uWVR9+YZUA9o7EBWMtcYquNLGa
BX9G/kVhR/a3lplQm/GMBhRkfhSyx0sOnKxYQDmnYNNr8EwE/p/79cbi4t9scR83MoAqjTvV//+a
kPlaIw04ApyLh6aeDGhdlhqqnpdK5ystRl5iJo6mTKqecHdIp7dBD6TX7UVICerbM+9ovwpXW1SR
WLMzBJQV0NI3+HjAy+N01++N7t/RlTTN6nfKsxph36EyhSXTn+AlTDWcJw6p9WGsAsmA3ikNilLu
W5NTeJsz3JW0A0zI4y5S8l88fVxOLFPTIw4uA04QJUkKL4M8y+TcJIJiyYCSmRVVu+MZ3EnTMdfZ
lsUVJ7OIS91WAZr+MHJnhsSGktqx2LiNsiTYXvEdEsIDu2z9oVqz9WeJwfu0l1avDiUBI0EBvtxK
Q/HsO1NXHeg7eF8kfLcp6pntAI5GbtLELVpcnpbtAZpL2D5TT5GWvUR+14VjK0ybCJrHs6Zt7RrA
uIRwKsEdL9dNSywx6Y5cz/4JRH5WK6TXSy4MhjwL+Kas+woWaCbpZTp5YmsJCeDchlxHpcb9eR2l
+M/wnS/VKH9Y9PQEurFXCi0ZhHqS4peQToUMh6EJsO12KBEj3JNWy2eGyI7w41vHS/mpjQL8Pul0
yeMJx3oMfscP3SV2d7ZgJKW4esyVTgfACTjc3gQ2xtxnVwlIMQfZGL0ul05wnZ7FQxzV9xmfgmJg
bk7F8wfw3Eb61fM4PpHYMNibdWAbh+m3liypu28FyDimE8EGYC1bcE+IGldU0g3qLvp/nLlCtnsZ
RLsMl9TM297i/Yk0hOffdYYjmKmr1Be+raJb7NFjMXOOb/0aPgsurfpDRup1yu//IdBr+tAE2p8J
Q3q8E3Gkq1UsIIWPc5ItavVcwDoWkKXE6dp151dqa/KaqCgpVnwbMjI8FMedlLxjws1zE0eoFGAA
Xr8TvfGW0QouMgqPMUCr3qw8ouxwXy4as+Lv4WNhsI5Nf4BTenvFCf6JTNjnq4xWpdb8SIOpDYOa
Y655H5OQTAYfByEDY6lg30j+yTv47SQVG9f2ZL/XR7wJpVeGrLVUNfSrjn8f4wOcZjBvXTWZOgGa
ArbuAd2MF+ACtRz3etD6nVjEdf+VWsFyPPd21N/VvR0K/AAnjEyvl/1fbUety90HVH1vZORk5YYr
v2jr3eoQfsocNLFCQdKCuPaFFiSGS9ezDSXMDXBKvzsKw5ddU2K2anwUauzOsV3qF4leBLkVw4WQ
K5Nf94DAQkDqzrmZBZ+3C2a9ry13oxm3I1aZcz9DNlLjSH09kkxxgFfSXmk+g8shxAHLOY1n6nj/
M+2xt34RluCRGcDMBrThQyxa9P9C3UT/l30ujjZLkNUVytm9CLIhkDKDgZANn28RmW+i2WuS7qQ+
E4psFNBm5/c96JusXLtJ/k6G33ZR1Es4Cx6lBpUdy5+LEToS1VBtHJQqwJCEbIo0pH/ggaa0x8AU
cGzC193Ko6jC1jMyuxp4CU3/jJ0fegN4WyOkfE9VGV3mJMuHRNLAa5RF4ssAhw04CJdRAU2dg1oJ
a5rFoURt5Kbi17E4vErllgHWYqhI+r1DfZdJSposs6SYusHGa5TpcqknbsFQYn4OGd1plDDDiaYY
4oENG7vPBEiWwQzgZsQ+oJySZ5D+WD7J7NB/rPST1I5zBG7ErU1wPIYrLijQLjH0QtFmHdcLXwCh
JxInPYJ0M0mulDyQBDX61ekhAstBxDfzRVg5nc5R/j4dFRMa6ck9DVN2D6WelagNMThdvaC1NAwX
lOHowMsuz6xoFNu843xyk/y0OKB4kH4VuwnZRududnC+MEAs4oRuAwdL7Ie2YimgRKOEUWQfUuK1
+Ag+h1Ge/gbL5VkRWJvr3al7v+FGTMAJlxn5NUynqk3b1KKclL/HNH0NrrRqjo5sOgzmwEK6o/e9
rfWD/WoDzPIfC1TxCKF/GzilKl+7BEvemdvYhZ7VVJWH2rrkOzITzNfwclKpZUlJlrRjQhEUW+tp
MD1iZHCmdR7TQqA1hDeaHjrdIsgWZ/dWEEgRKO5by1TQzrhMur3zgUGcO5EHgQjtIg6HNuJW/XBE
HoXEb2J79fzFELNyyV5bMPDtvbin/qfo2jIlzMMbo1M7duCgJ6lw0TeCRMudWP06z6/ysdZDVWbK
IAXYFlLh27Dm6ZgVIbGTy0E3XmqQXZNfeK+waTTlt5UAWeuVvswWKAglnlvyk5163/t2KF0iNIWo
cL3w2IludgxkWip+ifaHb/I909/wnaSGZ7qZXwAgR8EsAdJHyvmflsKobnd4ThFaJs8j7kqp7PuE
UUj30+8b5JgNCn/OYuCNIaQpQSWdZwOKWOqOnQiIflnFg619KOFVJuE+U/mVHWezIBSGAyIsRMkD
aZhwdIvOt1DYV2GabFLRZ6zIVAObvSj73Jbbq2CCF9cMXIOcEEMuz05vLiK3qMSaCUvH2saA5R4s
f+XHb8xPZaFASwqY2DBVqjJCozY0AalDWlgdm48GDfTwWzLyjsz18Ffs3hezZQ0NUtI/VfJIP79/
h2sbkSml6Q4dV4NosO3yoIU1reFRta22c9PT2ZhDmTpfc6HcQWVFO66LQ+z9dof3dWeAL7RcQi7r
SytTtWHJz1vlX2XaqaMubBZA77Rzwe991VjGJKPu7N7uGDmVwVQJh1G/BH/Y0uoqoD8huE6977I2
t0GYzbopxtDhrCtFWbQJdMMANBytCb9uyRPu57tjOVUPlqoqEs6OvU/zdnAt50YYFnGPfYNoxFMz
m65YIZW4rzcR5JshOaKmmYdLxPT8iyyhWRYMCcYcGB94ClmhR5KBM7Gi9qdnM5kWHxjBqpsqYrXS
RlST9Kw28hZcibiK3s00IJZ1M9LqRGiLg/bwDzI/kHYgUzbJF+elksh/+B7VP1YG77QEy+k+XDOI
oTz2cYSZutJ/C/ubOm5emRRtGWuGmSQkgJ2pffY8hs41ixieLH4waOTkRN44DSrMf/+u3D87LaZz
+SpnPpDQ7AVwoCZcYyOR7Tqcu5VpTfRoojPuka7KwX3JoAMU0uUc8DFSer8OI6su4cycwm2LE+IG
75zj8gMisnzsz2eIqQLVzuEtAv609hgvsGWLDi1Y6Udq1HILAASx1LYcG6PdVAsFVywPgE1VeiL/
h6t3ywLAWn3HHaXd2n+tmr4WX7MPAFyujbJsIY2wIGjpbY2ET+R0bbJP9CvxfqO7GnNDQ0ItAXm6
lkZrgFEGQuRB/FKxE8wC1IAhIyFDRF19ddDWcKPtC2sfkH7Ut1v3kcCLcodV8NPC3z6wzBSDHvSg
WMxdvohd58xD94J2/KvF7wUusfEERxuzSQwady2AJItJVdTAIvX0Xp8Y5n/6ZaI71CZOfl7NfXni
g82idnq2yjfRbnKF/mUhDNmmK88EWlZ/gO/YiVX+pQZDnAe7j5KM/ie9xKY/HtW+Hxd24/BWbJAa
fTTsQsGUNMw7cCczCxu+twaEqpVgSBciXz1swtmZG02v2hfKFBIHpSDq4RxOTjfnf/PR7VcYZOK7
7vS38a7lZsyhjgy8R0sYxzZB2Q5QDAJ6xtYV1s9XJfDxdyz/fuWRi9WvJBi4G/6lEQxc2QozyXKk
3M3L6RBFuRZ6Qfr9EIlTW5Ly3BTGiJ/gokCKoA+mH19/Gwrzhgs20GIMk0rOrV23P+IAlBcZsTYB
GenFLU1HxyeOE1tkwIto1aZ64GD2pSYtuc7X4GdU0chUoKDj/ZcbfjDmA4WNjP9p6e1300pdIxiL
U1TyXHkOCQJeq+gS78mwBZJ28Za9DjXt0unXx1hRe8Vzn8QGV8ay0/a9YqzKCW2AGKoQgDV7mlev
EO0PgArNJA/tT69zLnZmgGwebu633VZayJF2+dYhyTS1H0Op3hzazAKR1hthIgWC7OdMes6WgoKu
07beIInxBV+oDgoeMlS15bNfa70mODrVRUdq6Cwud6T5To+5XdAUbmPpNCbPEeQq/xjgUbue6pOO
NyPr8tn8rJjr6SIDeH9FwBvj+C6+vXKiL/Mntl74YTdoWw/9xhHdBS5lTirn12T+k+fx5k7PsE2M
YtYf8Y3w61D5LqGEHJmMGOtOlG83FrQGEr7R2ElD2sea8qEaGdIjEt6AJ3iR7TM9QHHYSqmknREW
z1sTFP36tTptt3kReX4K3RdEaQl2OjThGwTGzpwArhvs+vhKESrc3J58UO2n4F7lJWqBA4EGpkzW
nfDXJqtT6v+MNDAAj8MLFrE9+toFKeDxX6oOFFb31n4RNdNEF1aauGLDTPNV5BbCdeVI5Y2wmg3F
2p53zoe9ltyF+a8dt4Iz0woyG0cQncr+giS0eeGDDf5lCNB2FNQhyPyJj/0Nj1UopltGL78DOx9O
KwaM/FlmRjsqADj4EfnrlJ5tjcVNhaCalPmBb5vdMVBcOO7acPy9pMhNYj4AuDoOT02eGj1wt9b0
xAwYpwTa+MFyl4FCsFt9WpFoP6bEG7ZaWf5cd1VCbO6Cmw2zRoLPreL/j1OHyLESERcYGJy1u+Ok
mCA+0T6+UGQGXyR+RQkQc8YEUi6J1pIyytklV+p/s1yZViIKMJccQ/yjbH/Xv5/5hk8fMR9cw3t6
U14+0sNYHHPOW5cJLuoVjVQLW2p9Erk1NPIFdlPHnBbDq7XDJ7FvTAOhRHp3onxlGwtYwCyKKWt4
dgBLaw/qIVpsYgRYD/yWXgRM51eAn3TPC5NQbmCmuxqJgZtUXpI2ZQ+7kz3GUep/U9tjvjz+EzxB
GeaLuU/qLfUQwIquRedhDgUgRgA4j0y3WnzxdQy6sHJQfrIYvOSjKtqZFpgMOKjEpSws4SIzjcVN
xVZ7OJGdr+uQ//yh93WmNSE8WEhDkLRWwTqMzr5ndjgkRLy232J7K+l74mWT+hv4YRgrT8K8RHT2
84jCRsLT/Xyz+aMZAIBfBM/MOJFt/FCalF3JNlYnSkMR+ugQFVmTEl5s7AVel2DWFTiXYzXYQKiT
mpGNfFPw9UO78CzqzMJgvkQQeiQzcX6dVuAKty5qu2ePWEwP4+bYmNSapbMfJReL2EXnXV0o6bn7
465wGO+rSU21QQCbJlLb8SoA1bA4p2eiFxLTUGjK7MizEAkVaXbyDBHnLP86xxdOaG9k0Bj08zkx
8eMic98HhWFad/3QxxMvdRdu5NLw9N8ZNsN1moUzaUMGQmbYekpnplWHFdYwRfxBVgGSfsvR6z40
95MgjursJngmojv7xyOMdXP+BMcnaZnec6uYOK6j3Pkg8lvK92IXb37wj/6oklQUgaUbjUQJOcre
z0YXJc+dYAC4uenyT3iLEXZUuzHDnGsJb3HzWAflGYpazYmfNa8i68TVPPYR0N38MKrsj3NOFrsJ
b6xXhTLyk7758Td5YByMsZCTZgHQkWMPNspPk42+mf1hezFUIR4JOjc1B3PiLoCgGqoC54jDQuHo
gSwux6ULPZ/qDJsSsByp2+A32klHx0hOncjfjYlOlGgm7auZE/jZHANohLSC9qFnQTCL2s54CU/G
1QhIAKXVQ3irxyNPTI7Mdn73EYbFJP9Rb1ydzYxpYH5ipkzn85mhyVAsCrSv1ITb+SctaTVtrtXN
o32eE52ORlRuIG+exKXY0/6ldRAAFExMK2kczAGFidVV9GGb5gSBXuFzyunMyUBH13DIdSEkkwiC
3oHs5wgcHz6vxhDogyCnVFFhtLEWfFWZUC3b2r/D5++rNJDMNeoenyCOLEHQ0jzaXq+ffa5ohN1s
mliWQbncd/HgVo52rud1IpIt4NhN2lvIOk/90UBv2jzw6Vxt4GqWrroC9RCi2fO8o5UEehpUD3Lw
SwOqVHo4/yGCWHdw9mbk+j+mAjIZ0wgJJLEEWAuYFYc9l/idPTYCxXYI7bFIv9+gacy76Z2b6C84
2Fq0EPyjwCLxBBezRAKb3of0qOpINJv/myyCYJPcWsMP6RGWLLeaPvfARZ7OquYn4Bf/pUCX25Vj
xAtsoY5DdVDyxuHxZikbjjcGl+Ylyw0+wHSqzEC0GoHftWO2P3kfoNvgzWOduArrtl2xA17PsBGK
qxj31ZxcReoXJoFDD02VTv4NF4FQR3wFCwe4i3tbVIuIFDLdTsuB19D+h1wOrlRc7iv/kYHloBtm
8Yy5sixid9Vf55lgjiDrS8VaBlPKtcp3NFOc2ndg88JtkceChZWKHN0lKDdWiBdD9BJ6RW3IlTva
RocBIM26mjr5NLnDKl52loQnwfGRgObLqqIOyObbTGsfrw96FRlfNjpEoJWofraVE1rLd0Tqqzka
AbcJDlAfXpO1v8nWcnJFJ215d0XawUzKlVI8HZnCNhyQ6nED4h8E8B7KD8SD5+eIjMYH1f2+E4AQ
UJA5dQR5hkC3iyyi5bor0z+VqZf7fBW9i27EVhmRUUKAUyvbpthUFmCP+TMAhxm+HUdkH0+46bkd
FH96KoWt2lDHuCBp7zGn2OeNdCUpvAFEV/OWegm7toey6Aykyu2TvtC3EDGhynP//bBNIP1St2c0
v3KzBaO/ZEvZlVX6rTMSbpPFkfkom4hJNP8TPFTtZepvGAeFgOQbrDxJRTQwyLdHzD2NXrtV740t
jiWrrByF9mN4e0OodPAs3LFRPUjLwZYhey7t7Qaqw2fhUWcUaUPRL+o3zIBRqpCXlTjqG5iDMvbi
koCPFdc2IAaPQSO5gnp838xW4NGzxjinbEOGV5HQ/kc1C2uvyZaZaOzDpGTWuu6A06FfKM+ejqzl
vDxlzRRg9kA3QLfmtP7nHAKS/iKvZ3JtWHVUxhYux78gyUgFbX6RLjawJ2dzMqnif67baZV8GZSE
1o4RNly7RJrqOAJNfCIb1FZxvMn1Kz01Nxs/t3B/m10++5HiLG2ytp8dFaW5wpnpp7apJYqFVDov
kTUyZq6CL4qxwt8NcahY/V1dvYFIkDVJkP5QxeVfTYXHFLnAWQrcwfq4lQV3ixoteGEEsNbrqX71
1vNenI8pWndALK1MZ+YFs8IWPm4Mkd+jdHOVqcUs6OFVooBnX7Z/LO4G8VfkRqkLftWIO+OPiZZj
dRG0Vf37wCLlzaAIT1VdCw2FD+ZZA/FyLXampPzpzf+1pU5SuV94DeE6Ccp4yrH1u6AKpoyV5Rcz
70qvmVuKjYHxcLFsxq+EHv+uZTW1UId9+5yrp44HEDVu5St3Rj4sJDHvbRfNSWxkSEgNWjUgON1W
qh9LUk+TRpOEbdeSZdFePadV/l2eveh6524XUqEpw8lPbSLizcPegGY789ErFxh20qpDauwEdtdw
le+XUdqLAhV91vDiOYV9v7GNxMUOIs3SKzmX2soRb+jV6rOPybrRureO4lIyBluPFxvqXMjNQy50
bGVoR9CxW4buX+8KdeOAXmJBDXmguY3npyvPz5S+6+kLVducmQxzorxZaFWh4kYI9LmEcNQR5Xlt
N+p1jHxsB3JtOLBqYKP7BeF54gGES8RdM3iyy5pD2hIhxbnL51dUs66RbdmD7qnIWu/jUneXk8x7
OIrDA5MxkMrtSXF41YDLBeux7ilVzip1x11PcXfdbaortNghYMXLrqbNDts20gXyqBsN9zoq7/yS
FLIAqI2uf4ct1+aYjiSNYleU6/CT4K2ioljy0zq38kSFCCeUHzktW0zBDZVSVu7MFZGplCxcDeZm
JCO1FSm4ez9L7Nocq8mMN+xsgCWuOMUqX4iE4gAMtw3HQIzQMkFEB4uPVfkEhBsgbmK+CJ5bhiez
ar9D9wCBXDAZfoEOFdOZ58n/PN3Xvc0csRStSUMtte3mF7pYD1oo1xPf8W3Dk6Ws/Bl3PtMyEoPT
2v6Sa1+hdYCf2zprhXSgqybWtm0UM7yQgdW6JEJCigXIL4/B/TjyKHsJ+NEwxUh3eW4dR9H30A8b
DCRvcor1Pehsew62ewIluBDyZFLkLrLZUi+dyC2srWUjN/MlIRa7xW6J/kK27h62NGKb1HgxCsYJ
d2Vk85SbYmJE7E5+AvefCjO8lVZbNflG1A5K8C2bhKMvte8fwtkN64j2F1+qlsRjGPkJPmxzDP6M
CjNC4VgREUgrqgRrOkIGMZltKWrmWLcHfjNRCjvXWgWGh20mkXO88+TUBZH6AeobGmWN/aoQZBGH
rlQ9JdpxD4je7zFON1+IzZjgKiyVJEmD58qVA+RyM1uyQ5Rxs9WkaOW7w9UE0g3mbhLddkQn3h2q
AkYIqK4+VceyxKMLBRQs4RNzsU40MBowIA08+8XRBbITmKZZdkmUUnyb/Ua8NgWnRid8GOSnpmKH
X6xNJp1FR1hExw3fxU7WPrlfv6TkWWrNPDxjdV7u/B2VONxz3ffZRaruSBI3JHfemPM6OI0kcVZt
hhkuzOR0iDsPiN2qox8GKMzYe1ZTKQvG8DmC1UDJLiG5BUz6W0UyKPwpl26EmeQlE0Yc+wqhKRsT
hv99DTmlcUZS46ij1MiPCEg5pNvQo0p+/9/36xdckwgESm5nhNOEkAW+l0yOI1qHsW5Ux71eylcy
u8Ckf4Z7vFviRZAjAfvR1h9aht+XqoNHyEG/hwfk4LSBdeMOr0EjwXbCsC4FuUFNyxv6ei1yxQho
RXvhIdeuFKJEvQKyM5XzGkL6XEsDdld3DDIhTOXeC/x/hLDLfEYFkgmMx3VW9ELUJOlqr3JUj2uR
4fASaYc0oVrqglZBnQbeqHPVtLiralq/y2S3y2HTgg8NTUFaCz3GmDUkepwr+6V5mNo3grtL6j1a
61kOdW4oTdUeBBSWCBuGAx0cekGupC1PT7dijJrztrtFVvO57uqAyPnieRkVIpF6psc1J6eig/A6
c9CK5b8ASINRs84PViHSEdV7w9bDIyk86a3NgCdXfMnL7phhHth5SInq9msHKb+ob2kNhVTQxW1S
/vgYSJNUBRfASSePGstzhOu0Oucgd2P4YOrV0iNOsn08bUOCh2ayefRBYsLg/zmxUi+p452/kOHQ
3crG7Dh3IRPfp0T0IvzntLMO+x/Muv/JJZparuXD6FtD+fC9SFYKIWZK7/d3meAGnR+UwE4s21Br
WSQvBpe0yuHzqT006qHXzTtjKFHsy4BaThP7hx1231EMcnIY1OoDxXBEIgb/P3wo0MQjna9ZnTJ8
gYdTWTQj3m2RdF+4Tq3a7IXNBduBmHqkSa1mh/RKg7j2+kF17ECR1dcRdnKdbypGBDTFNQY7WqQZ
lWKp8PbXOwJlGFk2B8Iywihi7FXbpcMwumxT6RRB/bLXtU2CAL4nFRVDLraVZ/bAfXZ7IDxzO9I5
kyfkd9guhaiz3p934ufBIeiKNDfra+ePGqWk0r/VFrRwfmaHPVqH8/cOeSHIx6btAiGNJW6jwo5D
NzpLnKuftWtgzSmDmrtbmHJkHUuvT2WRydnGF/82jgKbNg/Z1h1iH9+aD0nIpNPc+FVst/7C0KZW
eku1XsJ1b22tVPRziS9otY/tcDaSl+skFjGVBGf/SkFlJ87N4lRWn2spGliOSZFPpY2NfeT2PTYp
MsVlMoJXt7jgAKoYbhe8XZZ6BxQhW2T1aFWED5x3dq+u2u1x3NEAobyzrQiBrb8f6OLc8p13NGPV
ARfLeYCb3y7DkYpIhKsaOUy5NGlxnWHX4NwtzEUVxKS8bpQ7PtQOEl+GuhfNzxBa06SehTh2i5P4
foOgQu8ILJBh0+WXf+yCtsobajsl3N5+e9FtlleR1WvxDPvQ56eOzs33Icgu45yx9w804TS2vCrX
++CsrnS21gzYR3xELSKLMKqUijPm4Q99TuN21g4sIcsyDSAivV7bkOQ0NWZs9uFW2GFrC52lT5S+
93pcCp59eI7zd3mP/INw5lL/ocnoGWX2qvJxJxbfzlSgiR4Xw9z4i81i8B0vbITnfhFzS394ROcA
fQVe6RoBpjBKjET9aD5jpcYX6EyPKWknDZJLrInRQBvvJL7YQj88PcKYC7d8Doua8cHvTngVszvO
PZ/RzcsSf/eDnTIhxShaPiqQF8EaJVC6mslqMTCK6dl6nyE9w6AHjiKEUz7lz/z4poTMzOsc7Brn
W2IYPpq5n+eFzLCMYe4+uGCywa3csMRhxzU7BNGIKuwRZ4Gm4N2tmp5+ev/Gc9HOcCRzZsOhJShk
dIOmw7AEBqOgHRvf3kL1xkQmJ448+7c7atAiIkRlQp8Jae03dzs3px8lzk0zLebklSAOiHLhz7qU
sjag9eMCBFgu+wHdoei3TPkDWNSxQ6fFuXCdzaCcy0qhBq0oAIwsOI1pPYvKt6Nokg37522RBdcm
JoWxAcAl/vwXY55AzmDbvQUZc8UdX0ogRyTht51fryPJDU4MsG5L2944taXaHGg56H3lm5DZYxOj
PhhAyFl7aHHx6/79a+pOGegOaMa2nB+j1Isl0sSno2O9h8xAd02jvRpPp+hgQ8nMLp8Y0kD4Tmrb
og04wkq/NahipMQ7EzaeFhcj1e2ngC4UqLbQxttIb3H83W3LgQv/UbwuuS7ixkyx7QKUGAdB+JDc
gAEWLM2ZD4Gyn3Tkdy2Rmdu3qzTVNJ3Ttb+0o6C0a1TseWpkBkwWuFh86Kve70oN/agYwd8nA/kI
9rSPUBUdVNstwYTShpEIy5NpugIAMbHIIvliixkrYJtHLLeP9y6W/5QdHnd6JnrNeg62jZEHrtrA
z17t1k+3clhuUP8OUCc1xMz5QPt02fFj+0enEAMW01D6I9qhGu+/iJYTqdcnxTqpByhveRhnQOyh
jsqSZy8AkGVic6uTJYmYW86d7AMrLN3sdo/j3w2Sh/r8Brucr3mh0WXtlwGhnhCFNAMxmC64KK59
0YmE45z/96UDboptx/51vXCq9K836Q1eFuR4Ct3piKvFPXeueEMlCpOytosTXM7oW+Xc5EqH+kI+
OSm6zuScUv7LlygPnhNpA8mfBRmIZh5OnCV+QDGvX9xcBXukhWyK665a/D8imI2NtEpYSIbfs+5u
ISJL/ICJjaNxSROxBeTorjGwMqC4evnoS0WxuLMhLdkhNqprJ/yUDDad5A3gIhvrigso+J4fivW2
dt5FqJz+aVt9nzhGcIOEHlSFZKGrMwtIxPpVFwARoMz6RS4s9EyFmEwa4pLs8QdCcABUjGmbQqj/
EOsH1WfJXMesq7vaCGm+4GAUcKd6ja/P+QxLaUcg9idiD6Blty3N01zhyvQq4/ByXFmvOl0wkDv+
Fhjz1t+5AINoxgtPxRbEQQvuSgHphDzmGaKZl37A7RcW6Z+7SSVkNKRhO72uXoYcZW761UElhFNH
cElBDDlyolRbbpAyCnzLRORH7mQ1s/fjYuXLyrs8y6q+n3S7Kh/4N5KTTrOrJie8+K5lqZuWYUMx
LZ8xIApelrK9vpDp79MH7U4qnvB5o8n67er+Yv/8pq2jJPC4yGcGz2aA4x4Pu5Fl8l70avMogY9L
sgjQB9iqLOv+/Lt1yDygRr0/YFPu3ZvwmyuKg38TIiyjpm4yquXGfseo3H8udNwWD2S+Lq5km2CT
+Wu9z6ZFCxw0NctMvNQGJpaHs4H1ZxJLmOV/IKrtkX+48WatuynTwN4d7LqhJ0v7UbIfN+QfoqFp
zUu1kJ6X80K+o5owtl+0LMBltznAxq1yPMbvCsx3089ImI1yq6fzkfGzfrsyknrLVQzlf+tNRuzM
ALm4578Qg3jdsWrC9iAgTsaXUvYhkAWY4XWJbXxrTyYczFA5lRffO7I3vY8MWwa8YwR8o0aXn+4B
FEvS7BD+Z6eebo2ezRFj0EejeKMyp3LouUQ5o7/xhobwbfw0mxZeVknexN+hkpEif/8OpN2FvxQz
4V86FSyOpANZhVV4Aky65Jed8l7lhnovZYyxA03/8+GOO5niCid5bL7CmoTKqxs7QL8jOMgqtYib
bFHeYnnjXa8J8AZLwm6wejeRtY4pE4ENGNdMb6KKhquUdAh4o+IliJREqO5b7r0OCvm5x+o9ktN7
v5QNdQcVAj+n16GYJPbB6VePhmgrejf1S/nmadipAax1+CU5TRKHclK0O0IKYCz3pIIreVInAxlD
Ur29EhzLVKLRTIRsdUAL3a1e94e7lw6CKaClBd+C0w4ToSxbXWMAFH4dfk1e9WlY9FcpgyQ07zM4
rqrWq7/u1RLAVEnaTLU2WvAmt/H4CLyYbrTZzCG+sC87C0++4yJEo5kFxldRyIGT//ICq57zchmD
uBJ8oB3/j/8m/wGAm5pTvqSOklrYPb7zdMj2dlQ80iYhSdDmXB9oV6QdxAj5RStI3aFzcOBCTeRN
pXcDjDQKn6i8dMf+G1mSY14AKYqtoes+31EiA9d70STiyMhc7DqbqLqAy6oPpTgN4gGFCg2GDXJE
Fs9XDHGyrNFdyzXLEU0PcNBV9pZ+0dXUACRLczsWg8Vj3lmcomrH/41BEz49n3GXBWuJTM6kX5IB
MjKu0gH4sbYv8260vUkbAAqGE9JqNh2Oxedup1jMm+Qjag1duJ1jnmbPXjEYCcFocb0d/nDIaUnC
Y6GVkkPY71zF8fI+EUUsCysBezIuIBQsNWXZtO5DzUOFT4olcZcaomNi5KRXAzsQ8B1DfqLKm8ET
Bs1Amau2i6vFlX7Ic+FjkozcVd1I63OLnx0hBroOjSSvyc/MF89AfT5yBeYSXaTvb50UfPxBuP4Z
MhMLmcm5CXLnjL6B9WCg7le+AMG+yBkCbJnQxIJbAxptHUmryOqBf23Fdl5Arjij5m6ypRlyMCbB
zaPT1zSewoOruAV9boSA4RQnEcL6LHqH6Rk89eiJav5L+UtktIu6xuLqTswSLwciBPXqet+8JBIX
W06N1/xhTARuNM5EZPDC1Q3F8QrI/QofkuE8ZG1KQAgEUBbcy/XghyRVno09M8GD9EvwbrEFoGVM
+zoLiaRlolPZ5p1AOhtGGiUtrftrrFV+F+6kyPL/WcaX0mMvCX5lnuwCG2zFszTItEQdSemuAqwi
ECdFO92PeR4vc6iVbHO18bZ9EyHGSz66OjlyUp+sjMyMOx4dClj+DCU2op1gdm45jga3ubX5j4Dn
G7NJ7sW3ELTCbrGjFzP3eikL0MPCL5KDwipWsc4KTCOlxonaC9rMMV+2pDn6EVizW3FL55YDlJT+
My7ruXDyuRtbPCx7a9xZ2WWVTSdMkutqtX/fXNUY0BuY7yvjSF6dEfgejvCmOGRV/X95fXMNUME9
5LOcrqpL3sfdC8Md6g4x1M5vS9WgegisS96lCmDgicEGr7vrihFnHirRw7qHWmgRIqJRjoguhmGO
YZk/QGkVxTTGFiIrSnYxwnFci1DoGMY7MBUa1gBu3XsTw7Y9v+xKHcBoCA3oR97gisu+kGEPnM8z
k7IZTY0uTQl1xhDXzf2sYetj0TLmOaSk1yBWarlS0ypl6ZI/IrqmwyKBuivogU1ldzsmrOVsrHK9
PfElj7bl9ahJoD2wyGUDw4vMbQ+Eav6FZtTMBN1V0uqg9awtM+n1dD6w5OAr7ahffX1saxDFR+fl
8ZGdaGPaLc+WFso2Xp8HaTrAPJ3IqGsnIs0BaWaWGPeQeLQSj2X9Q1cPKJYL4DiuFVL69tR1Caz2
O0oQ9KwJ8Ump4qwt9TffSboFZ+bTTqcKmxUi8n+TS/YaJG0TPBKWUOnJ38FxcqScoPFXDwn9r1HY
CuvxjZO03O1eSrlLj1j5/IeG6lJwIKJPl+fHkQzW8rC0r/BEsM1mu/cI/XmWYz4j93+kFKzSqag6
eaSp365pgDU3/65E9nwyIjV/w5dnyGr366ULWRFl3pUTVj0zROJK3K3dUCmxG4Gv2lOXJYh5bIgw
mbCk48vpuAKx/zl/m8vro7PuQUoet8MDvGgDuZI0DYCjeZr8IoTuySYvn+o2d7vdGBXPBznGJ3dC
tFhFC38BvLh//d1ncP4N5wIQIgrAXPBVD/bmJ/2Aj9OqHa/DJjJ0dLt30VHhnjFEzhz1BMPOkLA2
zWToWmK8VCNPdv2KS4jOcfo8i8M3N6u93nDC5vjSiXQCtM0gL479bsWMe6JtFbqcgUZ7yAUSMp2L
fG//tB3/2VGp9iW+FPg1V/HxI6H45JMw4EF8FtyNoyWj1KUAHowc6+0nq7FrWBQnYc/IOH/NSin7
Ffht0ATT2wdcA9xz6DoL7Ip1aGKkk2r9piIbtdmPaEhtV3YnrwBCYEUJpoRlisdWd+RCP2ejI6Nr
66GiNnEDpZhARe2dcPpnP6OjxQ52NFM4+hMYbjP8Fro03XZawMUYogrxwol20XLssyTUoBQQX0IS
8lw9rWSFPhNeWMJaTQ5CrYbMie6m+gT5Z6Ighx4DDtdohwHYnMg2T/ZAN2oMOiElbmc5OLAhZZkT
lWtFWrgmewp4ix1qp33FfXUQf6ITFgYc1DgSiuhNMW/R/Zv6Edg0BBoemJpc6fgrvNwl0IkZrHof
YhjdLmharkyozwUbeKxCYY20rDsZfnQUAvDf39ZoTBmY8sk4ftO6PVSvdgn6/tkeo/rmUQb7CiM/
a4vUtYj+KnztN7dfnEMHFPdkLr/g6H/dd3TGUumHm6oR9wLxx3P6xKAc27lO9cFTBpXXiyhBWLWd
11sBXHo/6S29lcU3bRLA5vOL4d4cZlZObR4uFWFEo3oXfXLtJJc98LiEeeLchH5P70DBri9oeR8K
TEG8IcP+f0iATiku+Fr9gUYmkG8gKfHcpq9IfUeOZROZyQjUS+lYdSVdHZdZdQNWMRecRnXR2wSG
SuVoU6zhyMje7ZlVQqx92Tr4ZTJaP+qKgLrqehE2dQAH+BPHs9AiWpkVSPxnE+Wd+lf57XqUtpOt
kSS+ceGVmXXOac7rkzJAbQIRUFvpRIxJwl72EsA8x2a8lnyrIDCNT4WEFDr+2mM1Jp5lKMMNaKuk
LwAOzYpnKybcYrd0I2eKjqEQr23r2sIFJgY4BuAUdJ6YYYgoZcu/gVncDW2KLH2r5jAt4z0kfOS5
3VQHP86Lbx1R3dv92FpLxxG8GQyDQjoglxxW5FYK4yRykrHduajxnw/4uOdRMcsDGM1Rw51oxt7B
s5ZPAiMhJQgg6eiu0/Yv9Ek2BgO81XXnxmzHE9zCXvNumyXQ8R+O15n3it7pAMccPgzFtgu0ryD4
s6yie5RRxs1p/vJqhicnBMgA5MrWBXJ5ZWS6ZNujUWh8fuTSuV1bvj6Ua0zG4kJwqT8BrKV7o6vT
G5vV6DfXoTx1LnxsC4/CB/vKzEqJFMAM7WT85RaCeT/ZJ/goP+QCwaAKNyodNaDD3df+fNCVCeI7
3f6ET+WD8f/Yri2BSYYXpupki7JMYKbqbCZqcnz95n5l05CGceyBAmJOQqxGgc7H0lh6meANoYmf
knpWTYXb2tsSY9sUyOzUXWkr7RrjtKWpDlT3Iev2nQbpogNL+vRgndH9+uLQ5Kja9xvdMYnR9yFb
6zyFfRai0p8Qpia50sjm7uYKMRL9D1Jy7cFIz6p5C0RjCvltS23yyKRCsQXa+TrKQXOZpxQPUOaI
HTn580GvoksqdnhQzi5dcClzc/yRssLb7WYBP/3THYmUizDhJUGrbzfmQ+Dm2HORrRr77A6jBVBB
lkfTtulCDEs6uV2oZG9p5RGgXgpw7v69lFzAMl89p4bP3UG5Sj73JGZWvRxnxHEOHvwWJ9c8QC0T
isZbcDHemXVc4+8seTyDg7LjVFOt4WwlV3qYDKPikoJUYFZ133yfP1dZfK38oeLcjOVIF3NJ0MTi
SKDlYI5wx/TDTfhMnhcTxscTsUtYMNvKcho0ODsYDuXIyO2yR7JjznW5QxDMlZj4KiHUF7X2J6u3
gIQ0ML2Ujfdr5yx6qULAsH6lriU8M7TnPbNLGTwHUHIR0dndT+gyACsgeH0sNLChHqrkffJ6kf4T
3EfM8oT/hJnWJC52LuQ+FpP9lclqX6nsJXjeQxY5zYuqWxbSLBfqxhsNJLj+aZikxt9jDqevSMPW
as+Oq3fe+zJV2Px+8q5Ap7jFHf0x14+WiVLZm2McILTX/NHpRTcPqvqwa4fGKKSelM3Gmx/QgIRR
+diLp9Sdps/UfQ3HUlwjsYOitwk4uqLoTrIdJe7WUxqI0EeihrGOSkDfMTPdCCDcQ6YlwSLxw6kn
Er7VfSs2XvhY8Uv/9kdiRk9A/hD8LUfEk/ERsEyV8RBblfyO9i0vwF9Di2qUFgQ6drLqxJy37NHx
7FBlKuAxh+ka/0wff0WN1CA33Xmt0M07Dw3Mwy1NYTjSj+PSLZLQrtHQqkz45N9Ia5U6xqWN7QSB
X90OE7p+J0GVoTweoClcijS+lHIM5974E5054TMjRwdtgNG/VbK7JXtHYtfoM6ndmWC5sNf0qr5g
+P6fGVFJAwlNl+PtbTmXTtnkfP2a0c7si7ARgeqH6ePiTFRvCNc1lziYahh4zxjGLz1ws6UQEq8k
QtzNtNOpwanbjKfMc3pjbGMpeXopJSMfrPdkAtLafxF3jAG/qjbArTJKI4zsIgOV2rYzoDWo3Znm
4H/ZcOnn7n91T7GA+q7aQ1dBsTZwlrOatyDZNCbA8VFxOBIS3nD4uw9jbREUOGi/dCPEp6tMlWao
xkHOAK6cOarHld2dnZEM7rvM1tN5xFcj3uKM0J6g9TkIVSDi8lsCPQwtIYR0aNiQxk2ztLOvsQsX
CWP4kTfoyr8ecZzV1juaXhQyS+EXpoU4nIW5wRKo3rwXcRwwVP3h44met8aBOe4icYhDrjvGcoBs
A7Z/Ue9c/8up+hcZCnRLx+P2/yptGe7esjeuw+/dLmEIssRfPh/qTx9tjP7CasCoRrRQRF+ay48p
mVCz6OzD9lUcVet4pc4FU46EqOmDxUQWUAK5gdcQfA9aUENfYoXCsiHotJQA8/sSzle5D+GtHwC+
q1iECP7kFT0IGKgKQaJY/Cwqk2av5goO0FSlbtmIDCl2GECwFEpnxqK+qYoCa7nv0FOLEIRfdvkM
mSbJlP8urWgNIHy39Cosjev6aK+gdHsswfHf5SE9rcZ/fkKK/bmAcG9lTo2F7rmOt836zPP3vYAQ
A+kvdOVF21HJFlWmrjRQJF055KvqIJyVIZ/KFdgxlL0HGowvZfdtf4apk7iQa8yNfR+4i+4GNd4I
k7pLDjB/9wTZUv/6yUnAQ/96MsBDxMbOGQvfZuPXVcGgLrabhPtwzRMuhKN4d3iJxZrUvMbJcuq7
mjNPeOGrLivt7JEKcnLY7Iy9RrT3TTgPNQrNunSu+dVVXINNvvd0c1HSXrXwghfXYhmuPW3gnUJH
OlOG1yfbszcAbi1Tv9tDTFhExQ6I3hu0W3Py0n0IdMA+pu9wH47w9tgIcqX/xfVIzq4W6uthPKAv
5rKnIAxZH2yHJOUmSvbsLuQEOuZJEk6aK2YkmZrHckifkh/5OahwqTOTfHGyUp2GyakerZGy7/KU
0vN+dz55HotChhKD62q7vBmwEjLFI10GEeoMNBHQ6FAXJ6guZUmrn9NWiAQmeHcCfRsxPLxYJHCN
fIp0fNt75USiYCV/dMi9I7MENCQ30xWnhLTaBPILALsQwbD4S6i7ATGN6Jp7Fy02m+DuORMIWz/u
ugdEmHLgJMEgXxW/OxUGMSbJGo6EmqTCILsrMleO6sLDVyalk1bE20YHMZvP+LJ0JnbM9KSjp9dg
7KdFX3XOR3E8LeE1ywdZ9aKKEBeIFE4JPZeSKZjRyV1GvrX11y3/t2JxPtkVHCEiEcD6ES3Ws2TE
gGkzSneXDww5z2wzvilJx9VfIIeiWTvhupcriJJgjy9TGaj6Ln9mnGwfKJsWkva8nU7Nb3yJvBjX
GwyHskGbqBtdVhXpRFxrQ9/x/YS1WsUXcM2R5o+vSW1Co5F6yHTIzmb4IPACTsyVVl87i+guZlWp
Vt9KR4+nwxQ4krydypb4poHIEQaXSIwfaum130w5OjFjb7maHGV/3+XTUwPoeKa5sL3Mv5AFe4Gc
BABAq2YEKHtXk9u8OpirB92eNCUQsoQbJFwaYmHxl2fu4H+SLpX0ttEjbOVveHhU/4CAFDI4T//h
CztubxIjUm62KfVHb6K2x8TfGHfKrnxf+Em5ZaeVG/PBsc2jiXYBDIuiJaeeohTCKmEQ7LqFvXxU
2y3gnYLaGI0I483WkcSz6ZKykkc7yEPAjPWnZfVZiezFe5aVKMaCIjqeTmImH6ze8hOCrv4I/N7B
di/0jEWReqrrCvNIWJpxDVyPEy+50aHPMRfu0qHYiB6PUE+xPshZveGYb/nzspgIkbImKtKJCLvj
+N/o0goKbnFtxQlCwszJadsz2QmZbyT+7lIs8++cclaN1lUn9PFWgKkYX2d9sBfbVv+jbFe4+BK/
68GIR1d6f3aWc7h87axFfmIs2dy5tVA6tVniOwkABsEULXtsXt0X1S1wGEtyG4lHdwSaYmdy3iTP
sDa/TEyQZ/gar+h7alBV+9P+6nlPhBZMRUBR8QoRsga7HssicwKLO7enLF09Z70Ub7m+msuaTTxv
+UWtUb6Kbn917XJZpEVDSV5SxoHrmKKwSmU24vaoeOrLP0zknrouxrwAStfT9hAOO5FFNfOzkl16
S9qfthGt4zgJTCeOWIdlI8LYsnkGenIgHuUW8JbqdAdClRh4dbNpDRvK1Qn62vgQBHb4TwqfocTb
j2oW7luLAr1dDU/E2rY57qjrWYbG99K2hT1/MPJSwZ2dFy1MLF1tE1+ViNACZ3klKxauNXlQRqND
1q6osyj1vGKKy2JVfbzyb58C6Zwtruz1Y4yo0TGL5JldjhHQ0VBMy+G96ENIa5lFJA10htVvaVre
71Zo1ysZ32xn+c0ATtrKSPoQvDcypBXZn2Al+3t44ZsHskc2D4Khfu40Iv9nrz02PWipfwFhOeDs
ttKfUknDvOGKrRBVJbqscaJ0b6RSnD0q1Unl2aZ5itRlMm6iNl1F9j+vDFsDVGSi+yZdH3NRjHHR
OAM7flojyfMwpd6VZXZm2EyHs5089wOB3tEVxaDabxb1TAXUlRQeNi/h4+g2LoTzebtIA6Ukyuxy
LpFSOK8x0LYmSjQG75+TxyIf0YVUm6x9EyPLPvjAiwxGE6DP4hDraf38HWgBC8S1rXOApnOknkwl
dVxfE07j/geIyw4x4dJmCROJD2SsEK522j9tvCeJFqrG7773z6/IedId1cA9AIfO7p/tMpfQ7zLt
QAIlqbf62+pM6lgWU2gpX60PVo3BHZ1Xq6/rdqEWudAYz2joOxhNItfC1QfR11WaKveV6M3AZ2Y5
JxigaXf9lkPdY3wsFzLJDGc9jRcFnQ7AVjMxJ+G4TmG34CWCvvN6N/i3/v2k9ODWypT4BILEe9kl
ETM1ITOxwoCOaiYFDnvwmqk6PP/qpjGw3UDlf5kZlhOJ3e73ky/2DPh/6RVh2JBH8C3zOQ1EpzJB
h0XpMdeMxBffFpCLoNjwvAFG32PZHeCpKHnscliD9ntLBtQBCKY2JyzGMhHKYN9g75AHDEqOdvho
XbzbAoGW/aHR1JzTbqzPCKQKUGkmIA3zdKEkFEEgHIk4gb6eRfu/qr19PA6bB1MFVM8HzN6buCL8
znpANmVpt9Byr5uLar7e9QHMC2R6TQuqJmshMkolNDr6ypvZp+//0Fej9DvNBymI1PYX4Cc5js6e
MA1FFci8CilGMhGaxLsDGCfZvEFPwxH0VeIjFia1owS7pFijtan9DIPIQDTU1/5nc/S4t+1RhJ/g
f5LXQN5iBHtZ0ofuCCA/ac7ezMcI5pnp4m1e2E3kmqtcNb6LnQf9h3DC8+CybzOTxPKN2nfhaSBO
OUIsNI+2xoFufGm8V2RuJKi6SpyjffAo7/lUhILRNUpVk7OX1JWofcM8J3ZMeWF4/KVSW/eR0841
8zxPkmy8tWe14BhgsywoK0WGW77VxALLa9FccetThuCGN/vUsaQ8i5Sdutuaj9jVmJZ0xCBu4xxX
tY+GJ0+uCelUo0fEctg5ZufTL+KuLCXnrxpIMnRVFITXQAncmeaLhBBt2r0hYomN338sQ9mvHk0r
X1Nnsqogr/sdbVKqrGnlQaaXzARHhWRXD/6wphhFiLlGPfWpjqug0I+aXAreU9RJJxxROPLIO6fW
3nRKm4DCGCylf/2eAqlPkp0+OKq34WeXWxTs5u8kA/ilXD/oh/wPpwHtPz2UQbtSa/Pu7XCxkSYz
31EEfPVAbTNN+6Y0CTDl4c6Si8kXiKxTf5GibmJ4s+FKvTQK+twDcK4VsvLx77FXToOSOQ8AdTt+
L2Q5OGIWZ5IQSFVkUwugHeOk53FUJupsoD214FV8/9MqShg3gTJ/THHlDY0/2Tn6adO9/zn5SQGj
OJMallYyzoVfyr08hi9RMEKgr38aI8KtGyNK8pIKEHX/rgw3jETVAqxc5QuPJWHq+oT5tk8/npf5
mUwjfrepJ5XV/5CkFqRFE6jE5mJudfpr1dYcjhh6PTrH0Mq9Agcpa54DEWqt7hKKtfOE34YPY9CD
xXRuZB8Zv6dp0q4QNjgCsiCmC6qOHrujrXk+YyGuIsln8aE2vdEj70E3c3v0wS349LCvySGzKX00
Huzu0VKhzMj5jKwQB1hE6gnjHMw/sNJQ2jZc6kmxjsx+/ofPAjajaojdGyI+ie5/Y8+VwW+gI9Nh
krrhIfeaDwIUBAcLeMwrbIYFKVaQ1B2dVPejLxcympvUNWQpJcwu1b26j4Qdi3fTsBwqFWysvMxY
O1+HbsAvnmPjp7xo0XXFfZm8FlJxYGbzansAMypWM7q3FY4l8ZHLHO+DXWI6YhnnPy9cfkgD9h+4
3fSOBe45epggKWcJsfD/bJoNR6a1y1yLUgm56WvEtelF7TvJKaHjT0r6RMK1NAsA3ATOKZlxRJeU
vRrPozOF8qR39BsXR7GTNFZXOLTvQhE/pk9JM9BK5BgmYDdS/+LQLBRFTPsuxUZyVN+rngRDcDlO
cibbDpg7Y0PPhdymfIpvCInbhXzpBAjMz6oHNhWCEoWdsNZeMDJWZCOxPErOfjsetC8Y+F8gsjZ3
BVKySdlnRPSRD4BkcBXlMyuFU7+Bd5EMVtUhOPE8J5pz7VJD3DKRAAnazWjar0ODA3wrcled2ue4
ZRqzVczd98VVTD0ZYl4fcdaR1rQ3f4ouOWaASgpx8o6d0ZTEN8uDLf/tBBPemIgZ8KPB9doZ+YZ9
GiEduCEGzPKJMEOZWl7V3g9JiTeC4t/Sq+S5kTVc1WG8xmc+MaPt2j3e5CX+/qnfI9/LPlrldw0o
8lFyDcUFodVYR3cOoSlbX3qHVrzWDc5/UuigyMCKiOaOMqq+/iYZWDLsxuwUW1OgL/3aS9ASixnQ
Z60x8oCbIvIqd85+lnXBycop5pie2SylstRBKYVP209w2WVYJIvNPm6Cpeq8AHXWST80hHQoKU+t
9nJ9AaSvUXTxDMUK53KDtXkyVkMewWGX3ZFGYyzPNs4ropyN9F67UDLwvw57CQ8syykrmqMXL/W0
+6CtWOh8cjj41Hnt3I721mUoBXZ7L/dVRyu1wguRWpEyMPOA3xP0QUBZF0de19jiszf6v0dmqKqV
beDUzHjPXQy0c74FQIAXJ+XRfzoqcl8fBdJDIdsqvVyn7zotAxhCb+cBlbXVbhUuy3sT/8St+Ohe
6kjWPHI1ISNjO8TT8msxQtZvKK6n1Rh8kl7wxHXqH360hJlrun4BlbTlrDQDTETAcKJjQHD6Fhsk
+9yieQaTrRn/JSvu59MmfDKVtgEFB9Rqp6BPtT7SStcKZwKA5akh6EttD6yaZoUOi7OyIcsipFIn
uel3KbbvezSq2+Lk9U6+LqlghoByLes9CXOIvsPtBAnY4cpl6II+FW73Or3gvzhD8gNeZtjz/4bS
6rra+SeNTNtSy11GZFPuXgAqB/JbWWvohUqBZV0/vNwpmlUVvixdLeIzgx2zF/83WmoIflAzzpHa
njo+WGsbt7BonMNkNbOR8vrbxYYKbjVFXAg17orNbpKvV7IuGHHCJaEid7WsmJIii+vOaYFpYUWZ
9I3XIUL4+4Tm7MWkfGW5BLFZR/Klwj83X9rR2jOEqqFj1IgvlQuXeJRolUio+nAtpoUdmovigaWq
VLA2zbpzKs2C08nmdYPvd8N7r4VUwjOdky7ZPGHFKUdv5SpN6E+JY3QkZ5j3ZQ7taapOza0hmccE
40wAYWMIOYZupds2o90Vaxz70ZPB0h+RLKvyb4wCK2ZdEZevTXvbAKBBik3MGfX9ri0WbtTHL/SG
urPbtIN53ckB+UlamAoBhIaYVcrtH5brkLPqyv3VmV0S0pHdkyeZ++JJTb7KmopYifmdmbq2MAfW
XTeGtcr6rGZer/vvRmZIbif16THFcYfTU5sGH1DcaoixdB4bp3NnPOnM6xB9w1mQyHHhjKJz5s9V
IeiILb6FwZboUZ3TGdDJfwaqep2fIvgR9oCCgjMfezxMpMRg1DiELUkaGaXC5Wdymi1FBpp9M+Bi
vMOd3X6tFvEAPvPQc4x0BrqSXZkcAJTi1IBiO4tJRUuTj57bnvTeFXrhZFef6SHuLGNe3r7swYvV
mCIP4VNmpeoZLx+tOA3ikVOCX22z+QnD6s690rhflAs9Je25uTy/nzRsPNAp/zPMQKivuFdWgJYZ
jPg/a7NHFZSTQGC8KBLNgfhQ27VWgiskvNbr7XAx96/hPeoVD5qBLBUrPYmVFdzjNHm+69ulmv1D
mhk4hOcKhYDNpzh/yJIwsL3N9dJzxdH4N0+4LY3eXddA1ruKGuLEltBiygLkIc1moNk+Yxllnsef
4GHQ5IRv+NwfSNeFSCw9h4O9mjPh0yZ8+MTojNbGFxzZGqUBBf3kHldHy+7aNmI3iprIuLupYNmv
DKiBJVNxW9ayVz5E73xc4Aug0Koj9tuV+tqwR2WweCq7fqiGbBnz2n/nabEM8nvH/t5wPxx3BtyR
mTCqkQIM1NiokCoufrOoX6R1bTeBqf02OcYh1z9sKcaLif4HDV977jOiwhXLJ1ZtEIm6kOpN/FKy
cX3+R5hIfyTr1GUyT63qANni7208rrOEOUx/0AXYCE8txi4Y/YR+sG3V440ztddXwRCUr3ygkYOR
Ur5XV/mbfHBiAWiE6TuB9l+JnOMDH/z50d6Jt6Ome1u6EI5xZtlK0PK+TOoD7t+FdBPT0p8K4FK9
ranwjKCCO3d/7CGcksuncZ55+GEzn1Eg8thc+PIKd3Fn24eWmqu0DS2ye5vrCjCwscY2JFZ9TuBx
fVVsltxN1iwLgt2LIy0uYhRqjSJpQigdCnf+5F1JhDrTqXlF88ReGAEyV//9eFS49RawDCy3M65Q
dPOEeGh5UJbgWbkDaFcVpA0e4s80IP53PM8Is1Ivv7op0tzidq9rHjnbD0t44KYA51qRK1ugkj+7
rMhT5BDM3mBEExZ5irUpT3nqTPYFxvU6O5KTytddzimEOLY8Qjj+b+B8iFZe6U/+BMa4bTXlXk95
PFmzgykEYsU4y459GnZrPf5YzyZ0OzmCGAi94Oys6V+em5tXXy5+E1qMZ7zZR6WGflKjQmyfee3R
Hx7WRCjYeHNZIqR/4w3UrqGU/PTbACViAorp6HKNF7h/NFSyBSsoAxLcqd4AunlTIg9xKkli2Y5W
ebehd6uQeAMVGep2LGouO1UvY27rerXAnlnC/aA+DOp0tbRGd7DmqwMWGXpq5DDJHyCiH9QMgmap
DOFETeQwW9uvKaz6rRB1SxcvkqGSA5u4lQBLPAo+9kFxi0EY7NZrCEmgR9TOgomdKZzAzVjRszH1
LMPeluV6VJADxfqgBs7QTNoMYstxnwy2JSsxI98QTBJa8LmKYXIvAdzTaE4KtAN5PUaU+3J5yAL+
ryFUx8ckSUzUwkqgNMqc3PkoiH5RS60aKJYPYWnKPz6/2UH0Z5MnUw9xZ90KWlvjX9NH+2aR+QXF
8YIxIVZL/oCPt/qHJwJZ+JInKn1BKX3Dz7Ah1Vym/9IANWOh+kKbK7Ej21GrH0i7vxEb5Dfnbz9X
14lmLTYX7ZmoRZ8zlplTcMPJY8WfsbmYg6bZpt6HnonFpTb0u7q8GPh67XE/W6VzOvxkE0mibupO
4EMKM6dly+qWJASAkf51pfujMYQQ4jONDpWwn9OC5wLzNhqTdsZCPzsHakY8N6xyEifjl7jXglRy
3U1iZh3heF4PREQSA6GDtClLQiolt5J+jLTXzSso946agrErOqA6cyfnCYUm+KRuRnE3iwZwK9Ex
qKYKsdw6BKL9boJZZ5jExJujj1bDJbdwOFXejMFdgZ4vgZV5QOMPA0cD8vpTjrbdZIn0FlVaXVyi
ODxBf25JPvE0OQ0RIPcgG85zUslo5Ql1Vk5GqPJsprabVHWtqpp+20t2UzA+0C/B8gvx72WzKORn
ap+Ush3aPnsBlZaMVO8qk5VefJ/E+nIuF3fKJo9UTRsAC2VdRfhvCJe+pgylcaPdYo52b9UT+JSM
7GD6Fng0R8LQA0D0HmvsLF4mOjKAGLoioTaI6PGHXCvv1E/ylOF7q2OSoxUXf+bH9RD5Du6ApvAA
mfO1Fj1mJ58MjIq/c28Q84wc+UWlX/Jxiyb/E5p2XJr1F0bhcnnqbQ22PEhmmumITclEmmcMabCX
bh6TnRXOTHD5U8T/VAl3xKtznqakcHj5K14vxuiRE03oydSELDNCTDgRVxVB/6f3lM+CPfeVKp+3
5Hpi2n6DwSYYXAN2MjsjpVnGoxjmKKQ15bCpizfzJf8rj3Qa/8hlujHhMQhnHvOmQxpx1C1XkmVB
uhaiGQY5pO7V2KJiU80bLQ6ROeIA/22VxJPvpBpF+2BpmqxrvVa3ecQ2ElJa/ywmhzb6JPrNCl+m
6QzRxGkpO5PmZ8IXqp/Tpor61eOpViA24wjXXlK7gMWHTBCYI4eqVLtSvH585HzOb8baHXUVS9Yi
hloosCzD6Lyc06DiMHx8Ux9G8hcQK+Id+TyqPiqcOlkt1bMC8jGNow5ITJKJom7kMrxViFpWlmHw
R8Ebk/qPaGw1r39g/Mx4s8nGM0TwhdTmDWFSzCtIkEBvLFAQ73SD5UVGe7VYnzLdPyLG2g6fyruQ
O32uSRt0ewZqF//sZBkHmwNzYhd/1W1kS9+6U01wmZT4W1Yp7dpJldnXx+oq1HpaXQMSb2kEVWfD
6IQsWEJjxC4ytc0Z/YRW04/8NeaQeyfHp0KgICpohIGTAj23O6sy5d4DOoHm5Zhsauw5cjT4a37O
yIyK20h0g02UxZzJRpBqsh0R4Scfb/ymJhiyLPNsMjrvhKfxknhFbuhWkhf8x/D855n5KF4bhogF
uJJdC9LBiyTKyFLGjyUvQiaE7m2B5MLOy/5Vh/cz9+5avWV+pChD6sbSD1gVhDXuitnUTFA+oBz6
OWqttL8Dw/LEKjZCH8D83p+jmQLuxFenEB5OFquDp4ZPrCORfU17/CkUNOBDikeSYW6pRV9HKNGd
2Xs/7+UrQ2SHdMAft4p3x5+2exWyqL8x2kCMDhG5TzMm6ifznupvmgDVsXidggX7FTSqgKu/Za5V
k5Y8veZ604Ed6/3gsA0MoJELfKpXIuKn/USmpOzhJ8zbrB15smrWXAtfAyQBsBAfJuCqjXlpL02u
1IriesTLF+JRknIhTa08llDdvWDJeLJR4Abzh2tLt8oI7s0PTn0f2LAT+wafzl3c9aJ3FPXbxIgu
JreFUQcJMnnGnHthaA+NYWa7gow2j7FsO1sYhaX4Kqt6aAe6bDzfrk1F+LA44Rs5O/2T+BzlN7Bn
s6SgKdLPUv1JR44FLgY/z+U5/yVICe/BKfvTeFiClzhb764oOUeNgi/Z1oh/wdis0diJDdK1fZkD
saw1EzTysg7zFhre/nppMdqn6jxiFq1NM9r4/7uY0vWcIZivK2C0p315VN9O9BuBjRuFOUqHQ1zI
avGYZK0J/oE3vKSL5Tvch13toJ0+XE2F2Kh2qpFCSCsnsC2KUA31tcC9nEuv7iw2Dh9REnflaDaK
MzlHq7qsmJ5Nkc/q9irK1RpBBkvB3ZQ8WbPBZ274oNlFyfS9hRgtJt+FRyJ4mw8eh6szn8vC4YlI
aGpvDNuos5+XZoVe14TpxZkEry3mRcxZ1SS4kWiztT6uoS6IpB3Y4iAuHmAubc6jvpLwx1xLNrfr
h+gUTZCNBpUmpi5u9WWk9wJ3pA7JAvQ00GVlonoBmwnUg17Yb1Jn1ArurRny4HrTQbX/2Pk+inGE
vOWogm4huFOKzOq6NG6llVlfuOoqsYJchtRvNFHjnZ7FtwGx172JERui8Et3autkqP/zmOV3BL+5
SCCHB5JOGygCQouyKqAIQ04SoYrSUcs/aliYudhzO8dhr/IrjpCBcCReVmcv9iIf0V0iBLkj7AuM
f1trk+LAJeGKiM8ZLH5Gn0WRp7KV5oo+lQnVKXaQ5L+79EdOu62RL+Y/knbk31+A/F+Oa1C4iQ11
Cywg9K/Y+FY3GYlyc8suQ60WS3OtLulTwvpfW3zcfR9DI0ZP+dtpVE6g1GDTuH7f27tSg8aBvV3B
SMzYUEZrAuJ/ULHF+9tMM5n8ojECxB/hoZd03ZGJun/51gdw+L1H0cr0YgWaYG+MzjRrk1rhXo7G
v00v8pKPZxmV+jkMzw2tL4Hk+qCHBgePnKeX6ak/8gqites8FVcSxdliiafmokXQ8ZD0ZYVGfWxS
kNO8lGvquQfmr2nuWZ8cq7dtP1bTJOdKfOBjjD9YTPN7kiaOGXCiXGK2tjsYW7hqmft767y5bQLR
5pGhX8d/KdBOtWvdwsIPufwlgbsfzTCjiL8PvvP4vMCSEKyr+kksn4HnggDSwvSwdYuYOaaQMW8I
jptyRC6TITBSLweZqpC0f6GZjGUUhUFOiZx/eSUNJMPmzSGcncwdD0cZbxBjlyfJWyAsJuAz4+VA
XAr1wbJsX4Kf0F2hVxaaYoDpx7y1Trp44FaX+hXlZbR5HBADfUpjqYw52MSd0AGNPI4EREga4pA0
hO6WG0V7gLIW0iW7NGwYYMiYNN3o9/Fdo/Fz5vtOjO7z1zlfGYEjewIjsMkg+wYBPxJ0yhI6vvXp
TE9AdmrgSZgAfKq8L6I6HtTRJmmeQCimycqO9C7S4NOBolwLXzYZLs7FxuEENUhr6C5ABlbG7Bo2
lQiedg6xnIW5xZZGH4gqgxhNR9ON35qv4JY6LhHmJBzQaRZ955w/wL6jcdcEUQPfDYrLzofU/s9f
8r0+IxXixUJ8OoCojyV3ZS20JIekDC1C/NKXV8JSRgaC8CzO1+jKJ7Nkh2QWYCb9UdRJq4eF8Xpl
c2PntO3stZyGEH+1PgZPjR6v591mDggsnxCnha+apEhDnygkYBBZj3gUidd1VDTur/umG/EM6z46
EEdN9FVIzT+3qOnne2tgEdhpVUXulBsBA6htRE6+tDvuqmX2aq478EKRDMGTdCfERlSiqXdQJxby
7bBqUypQaHU4jqb+xuvHsmSXmu/WLnrQzlC66uqrNxbvro2J5ajNWvvC6QSxVe9RTonBNENcTCp2
MPuY2GKvVylB99OpaLfveRn00H30jBsBDTWB/+DhiKW3nEZ2k9ypPAwocZWHqx1VPP8ehNfWomOB
Lo392EVgr20PKZWG3Fll8JWA9YNnTxf8TkTV41+CZaNei6Z3eZqLUUQJ38/i1hQ3lAD9AHWDbOxe
zUDAO5kzTT/orgK5WjG48UE/9wYUVff52Ao/clRo8GjV1o/micbKxfFar8nWrJP4IBOS2VXRZxvp
aRjbAVAeFe3fIxjoUAqbHFY+rgc+7ib8RDJsn14NtfvEECJCUMUYHyqZQgQY7POuiI68U1c2Q8yR
98r1VFzPH1xyUT+t10wWQep+rAP8zWjW0KV5tatF9LOh7R3B+Iv21/ae/MvlguXdHTTF34+JQmju
V1aJCsLcqx6PA/ukVADOHkrV7QQ/Z9DNhop6Dtliv+Z9cIgNOzYYB40qP95C1oQ4YyRZNQOS3PA/
EcEmqoePtRjkAn6HJI8gI3BMLWDUC2FTKZNJU81CUCLTEf+KCjvOoyAIm4167sqQ7HkFHhnQuZWw
yRFvdtTI9k1qt+eXnqAo1SZb9Perv/2PwNqF0Km6FntDjioUlFZZSesnYFWX7ENSiNtpi76kAfyR
U5MlBXmbQ+PTc9R+60Qio+aw5DugwaYqzerzyJ4FF5z5coPP+b5D5PaNOFPUTcW8ZpJ5PrUI9XnN
uj67HcpRp/J4Y0gU1x2SAfxUkZyTp9PwNoIZmGi5dRUmL+bVhLlcGRGhT5kvTO4oX7qgjNhv8dX6
rhq2d2LfqdE4DnfxNVz9hmBamLC35eZk6v6o/s40jQGY5bANEmDz8zBBDSd4/RnZS5h4Hp1X7EJ5
zkhnqYGmYxbnhdPfmAPacFt+relhTqXs4pBFUKmfHPa+OOfF+X8SYgcUKgsTMsSjBrIfFwaGiWDt
t+srV6r2RsDAl2ltxRcmGmH2lxb1XrVu0T5BxjYadUm2v+slIhC6RiA0aQEy6QIwSZ+VyNnESRxC
HyNtbUUaqs6UxD3OjQqs16xbvst7/bF5tsulnY2lgUxEYqztyYWGFVW8vTXCgSQc0dn80Q2caTfh
/2m+tHSdAW87Ni9oFlhQ/yYdv4vg4LjNaandgUlm6XMwNeB5akUKPIDtyyk5WOjz/1XdExFMMDhE
fA4U+/Nuf8mZvnXK4LSafDYNp4sPd7Gd1avrIaHlmdZe1+W+bYhvEOorLxhv+PrexH8Z7EomvFFk
Gr564f02nRh9prdwBZ4yO296zk/9sOKTp85j6qVcvAgDofyQsQ87GBNtY+3vmzJ1pOBH8B+e3wEp
Y0VpjM7ULVsT07E6JFqSfjMa8gM6oq+WRYHyyKELelalJ2nB/8HfdhySuK2v80twCGEM3h6qoRzm
6X/40XJingI2boJdDU95FefxNPrakN/Zb9p8Fa9NQQ6rT8UdcIY3kIMEKgITr/slqCKyXpR/y+Au
JA9zf6vS6exLoYTgmM+SCyu9cGgUc/+LNXL+yyLsK9Mee0BBxSiSLU5s3L61XkOdWfTpwu19ci78
4hrHDZfeUOjJLLDbQUPF0e2fi1phPQ38FrrSx1eRkiYV52kxOtiyToVDfN5R6am3LHKNSfxYWtiW
NyA08tu+TMH34Xvs8x1Gh3f0zQRNXuU17e9tnYx5xtDcQ14Hzu+YhAFBDdzHYKMQGQaNz0kmkMdW
+iehXlihqLGfeJYDNF/UDo05WK95ByY81avhkRK3LmQk0aKh71Y91vfx8/y/wQ2TW6xi+jgOP6By
dO6Ntx8mRWMeDzB++8VgBQfz+1bOgRAW3wQikIks6vNKwQHiqmfsLoQ/9hCS+YZDRLP1dRHqAwM0
8uTiotEjX/vUWoKPE99hRx195gsK07TIWGQ5PZeJP9sYXNFipViLl3peuRs+FM93IXoAf28aBqaa
Qva3frw6KpQdMUlk+KdLY/0Ehlbb4WtA+CHqc01DHY7VieTM/Y3X55zykhjQGO70tdaMk9LIU3O1
yA/jsaDcWj68fxzNMJYziTbEZgUMBB1HUH4L2kfkAOKjU+OMGKcy+CPsNwejzQtY0T5SYEsFPtah
i3g05a4oxgx6kLjgzsUXRZKxA7Z8O3Pk/bx5EuOxgQpOOVEIWNUmRBptUz94UtGJLqKXO3FZ4mWf
cP0IgCLGeIKmYH6sURgzLXSLCnL5c080XxQ4+P0ZAT9dY8o0EYDPLzpmoREYGDz4aPNenI8CCcq+
gmM1YXov3xR1vH5nTsPRxhGigAuuOe3yIYYGoex1d3O9ErNxbK+kqYxWZ9Ixasayb94M4Iy2PbNU
Bhb1Mpprpsbb6wGhff9Z1t5wGTrTQGmzw5e1EwVrPMt/2eJkWUvXP54XtUgTP2TJYYtDXxulyv4I
UewIwU0Dr+lhA9RaJj4oAlDgIfQLIVGdbhhLkqBABEiFewx0NVofpS2txFtkX6zJdUbnAxT7QLrM
HU3JrEKv2IzfdiVswKKXCKr8PNixiq5xZO+VY9KnNHvBh2AqZasdzu74zhJmyPTpv8dCy3L9XBiC
fxqgwKQu55ZFDyGwRkImTGCptMpQncCNZ4pwyqjzU74IVqc9eH7A5gw3Phee5B8OCdbexOZktjJ/
LRW8JvHBA5gbct5CAOX5bHsbStxT7LxGHtTVgmsLOEFiy8yblNwInhr1RZ5x9pMIKRdftmICYnPS
p72xpAefVZ7DIdyDI7YB/VFbEzY5ozr10rLw2mQjxlfSohsQ1PfB0liFb2qAWXfwzFJzpiIxtg6i
ly3xAGyPjZY4QncI/2hLo3pJoKv7tUMfCvKRQV3USuUG5Dryc3v1/sgR9q7ob7sNUQ/os4GuIU+J
cwPHp6Cl4PqE9Q9l6ZPodaQokkKkSPbbS9BRoTcVeCBIRmLDGgGOwxzOQiXpa+fayLgq28K3Mmf7
oXuKjKrSOhS0S9XgIXeDq+ei7EWwog79ZCU4ypoKNs80YH9M5x0EGZretz3Fc+eVcoIgn+Um1sao
0HRMRFtTDTXBQdL5MlJ980OKivaNK1vMwAzt/yRfdMubgml70hQ+K+26kdFlVuOMHiKzlEUAWlvZ
mgBORPIx8l9LFLWq8ND9/CA7q2GwdKLSDXf72Iv5LqgO5io+PF0lpJhoPFCd/3BmtMiUwLb6Z5y0
2XqMhdQFnTi8Y8H1/OxnmeyoSSdOytdENzxsUIVoWmpe6MzaiCspZJoIhYsOO5y7RNdHV5HvLVMj
l2jjg/e+KWONESDUsUU0stfwDhQDqLiDNbdYRhi9i9OXXZSsKIQyOpms7iUA2y7zRJYeYn5La3m+
elclG3z+KUgvvJJ7tpVy8ydMouGLuRXnSU5X53STkXlvNDFg0AtUmHT8NKMM5d6XWjpPcu2brwR3
r98BJmVSyrYY0qraOLD8Q16pTaizOot0WwCOZsOY6iwQROZtQmyvqG0fDlRpqXE52/6JXocdKMp2
FIR5qDm7rRQXn7g7mmeCIPVjVD3WildQ2TxlNrbqodFvlqEgY8WX/hVMI3W6FkgWhmWOz9CtEsSY
uk11wS+/CFWESC2J1Ff7f8ylCdvr2MO8qcQCeqXgZNXGmq/uQVABR2wv+fSGEoxixkXenCd7ZozU
4SlMnbPz/T1q0YF8eBNoHx8JByVhyAOukHH2gfm8hO+yRSp2RP6ZVoNUpwmDMiHvKXWu4FMk1MJv
hNqx2uqjU8vCwoCJQX6USj3uNJY/8rVNG3h88fLwf1kb1WZsOaKzkl3bUR3AcNJD+uWxFGt7JOe4
mjBA4n80IeuIKWSNgi8uLtK+cdiwrkdYsOMuA+UdFWdtKwjAnhOyYo5B+UPQo/HwMHlQDgmFJkzR
Yz+d0IXafb40LcTejh1Ud4uaR8CpI7q/z+o4NshW/TBbl1RNjcWjsiRNttoeF+44QOGpsYMTQioT
m7OlDqgJoedJkCzYrRvmlQGPzy/snPHxiV3RHG9X9Qo4i9jAzhs1uBXugCQTOaqhtzLLksxbJAKd
9Ico5s1n96HRlT6XJ5ehlXT+iL5POJdTk1Q+pnh6pW8SuU87fOloXNo2Gm60HsFXnv1lZzJZhpW4
gPMuQvHst/qUE6wlkP+k6t5C38CSj5aCyliAQYDfWAuodPdOMV9eRlGQ3o/CcB3+HGrF8cdXr0I1
ULq8xERWgVjayeLdUY3cY44b5nm8p7XdplsnhnhhV/q0C+CLhJUHrdfmoQMXOYuaARY0XEF1V19q
Bv/ZbNr8BMI9d2P4Dy+aj1P+T24mWtj+3qr2FE+yuYDrM/uvunzwgo4xaAWRUYRah1urobMMbeWv
aAFSxS1R/8wT93U19TK/rS63n9RXvFDwNEDm9fWilccWfhrJaWD4jOmuNvFnt2Y1YjACIAnLRbVp
ZO++ABu3eyjV5ovv/avy1QkOZ7HCO5/yC11v4qLdbQy2Gsl72Oxhe8sYq9e69wAfBdFdK4F/I27l
mfxKrSgRh6zKaGN2QxkJ4IBbQSOo9EAlT8lND5ucWG7sc9al8TjUtDe8D/0VEuNNk5z3trw9VMaQ
4L5avNgo7dYzNkz3WmsUPR/+ZC7o/RUl3kK8f8rMT+SumTgu6v4IX0F7h65oHu7SQbxPHh9F6zDc
GOpiSDreVA9nwpIYnchKUT4kb/cm+OVwrUjWElJ0nXExlzfFSSt62kQ3Q3f2M4yQItxIBDp3zcT7
2jcLfdO9owbJGvUbVgQdVpAVDdwdFFERy7YtTSl8XfrYkBe80LNMwx2NVYrqK8O5P6wjLYq8tcza
YahZd7W7CVZkge4W8BshyFz+fL44WW8rP5yh9xtP5G/4lHHwiyTp82FzCZxTM9YD0uCSsXFyGGR7
RGqZjQ+22ql7XxRbh9+IOPvAKx9nBMP6xDNtkHcnRnUV5UalePWIpie+GLtihPOwGvnywy9jJvhW
iCMtYlQuGsIOHO4cHdiiZIQPZ4NN3ptqTMMZKRoKKHmVXXljXPoGwnBVx4eC13k0sNB4fGswKkWy
i7QmV+5ZXDAelHXiUXWXCWTTHiGcuQ42oQbDpTKEMc8RvG8NBTENPedYQ7QOo+Wxvp0WzfdzsV7i
B58dPBEEpklH37kXoiypHnCNOgh0kGFyJtUMBpLAWaQ69ROnE3kT/UpZGpaIiBVA+5Y5jogAFkxQ
rtrK0gYQRbo4QvfB4zqxfrxWqKV0+xxoM18KTlTUg9RJlgbO1AhPvNPJDAUEnC3j/1O1YjegX7Ey
UaTq3Au4kHQoDwxEb3YzBPNSnoSgvnQIJlOcKwGBds5WajRBA6G1RiQrWFO2/kuYT3PCthr10Zsu
UIMdVQ9o9skBS+cIxFMfMl2nbVA/O1ondhEOcxuMazX2I6xV97UGPyNBdfkYD/+FZz1GeKueIiF4
qu41r1Q+7d2tR0wu2/muqS6ngsQv7XO2YNfJnMiDDuw4J3iw9aHCcfeKRpfY5uviRnGTnIH1GXzQ
Cph2+B7KYMlGxz/jrYln53VX/d2e5hEpSAZA5Pvdq7emCK9QPqfsXhTp4owVdl7V0NtQHfGLYmii
Wmqe9Bk+nwzZxudbvGpEZvInDHYBPDx4VLV6N84nlkOBEo4YHOaJZ3OSOW7L91dkXHLShPZcWKQi
EU3pWdZNCFXmkh9OGQZJmWSZop+6ZFLe/llkINtMOUV8Cg8LFONSbF/nc7HNprXpbVU1UUxoUHJk
UjwCfMEonOoL4Xx25HQF4JcQaoc6m90QU9wPi9NFU107EAguoTFZvAo8V4/BoZC1ItLOrhKOs8yO
sAX4Et6vTMEpv8MVotz3xaqcVMAT/IY3yXhfghP8ZfOA+yvInO7Wt0LHB7HfI5AdmNH3ARlwaql1
3qI+0Vym2E8SY0x/unv7fAQ9ZH8jwLtV5pUxhEF7QOREqoXAMFGQ3vc4i4S3bTyqsEVCFtEnaaDm
VkZD+zaTsVDsf9kbuDx7kSpR7O4mb16p2aBuhb+SdSe08aKNpPcW83PO4w14V2nqcIbuF9+rcM9g
pgI5O40XuZufVAjD55HXzQKT1qXKPgrGhjNpaU+a0gi2H0jfTLXOsCRmbTMXvXNfWMdh2Cp8ZSV9
rge2S0JjNlt1Ent3L9wI47PnXgMIPn+ErjPGABCihVzOWOu/pQfywzXXYKS6G8GYXnBnU7dhYOVM
h2mgdlDKaljOtr69I1VbZ6Fc/UVCzDbsQ5f+hqfke7Ehm9XdFfm8TJmxkCe1098C5sPYyVuDL3qe
b5wUXiBzZxwokmGfaWLn3z+b3bMje1n09TUsXg5rue2JybflsGXe6BiOQ7Pv+XbjalqVw9dR6sIV
6LkkeCg6hLNfNQwDeBuqxheSmjWwBvUJi8Gc035CGJ6QjRMHCxGtGj02N54LOBu4H4Br4K6QmXIz
VhXU39qpmCLF1nRbjlQz1Rc2JooaTgIE6hraPoENrlAgwjM1XzhryFqYuLy9C5mOXeB7u7IdGq/Q
PWaW43laqRoZCa+s4I6bMe25OxVTvNLI5UZtnuGWA8Ekv7H1B6T+TdREtWWbfFCCmgkZQ1iVsvsk
DSvRJA30esuci/12nxXBlZBEs+y50VRZLMTcRO7YJafr0ixp/D+hmOmt4QqYPZk2lgpfeuBOA7lB
4t0crYupdnNyjUUsrCoa7gj+eapU6wftQItrKSRqCz0h7Axqz80v/IPddQsSORA+9P9PqzJ02OYi
FxRXfaUrDh5YjcHXw62uhwnoupIZqObCqkS/LJXkH7txfxLMUrrxl+lNyzQHuebYCZ7hcoteou9I
hOoxRMk++qDbeHkpcTiuVKlOY0x7AlOWfHwIk20gj4f82h5aMNMaudmq1NxzQvNTWGR+1swdXDrV
ti+YXDhPVlSO6PEcABOoud2WaeTiO//3Hl+NsDwVdmYr8b5OptLpnYLX0GnV6+PO4Kb03s3P/3hT
H4kx/VGD7D69zVqE9GlnFR8YmDAD71hBjtGgisX/dFHKYEInn2fTg8W0Ukqq6bPWsxpDAdGh8Yht
ccHD2uzu8ns/JpQ2lXaO37O+2jTH+ud0iO+pzr/m02Twaege0UHgUoYgmiYckJYU7q19sIup9hLh
X2u6PyTU3sso9xot7VA3fxlXkSSpX5OTGNf/9+Pj3Vc7KPnv0ccqUKQSrTN7QwwwvE1htOh0B5by
z/8wtaSyM2GysPYM5gCEzO+3hSkE59+SuuFSv7WtyMBAYzrSjo70L8SI2NJ/ngoez5cWlytaGxMO
xP3DUg2ZTMMl6xAWixjaaRkrzWO0kLlu7t+V44hcphhOPDIOraYoKp87V0Flxo9pa0eket78WERM
zL5jDUlRm1D4N+MfYaT8+zNvJdRXX2izMS2dgHSDxq3g6wdqJ2bBPWj+gG3A9n+S/cUes8mNWCR/
lz1+t2iOOk7NyfltApIg8HM/V/NY4lHypbn7sHYazUU0RpMOCEMQ9uxqtUAjfRXF6hOhD9silCCU
+CvLw4hLpqEO8CGOMbI/d95+05zq+G1jB6ZnCpivHtWZrSiW0viAuYzZofBuvRI+aXC6FjMOCY0a
GIdiRoysFu/lcmaqCRj051SUUo95dBXrvTNtw7VFDXArEtseu4HmxOPXXSS4ttxat9pqThaKBB47
Fx02EvhFAbQDH5RFhi1N/KzVUK6ZY4Ab6Lv8JNUFty7cfYQk7rZI3oGTIsz6kqAoyYxjAVD25kmy
w2dhwArUvu+lhRH/CFYzOYw5ZXciutRt/+rQQJw/ypK9HsOOu8JtWZxVHLhHGS7FQJtIf1e7SEiJ
STHfmu/amgfOWC07BJ/VAvybFZFSr1LLhye5gupMbL3r8P1lgXB+aDI+h7HfBR40BiRJ3BpDUSa4
WkjIbaBI0AxB+VcahWXVNfEsxBc5Gy/cQEqbmnYdaa3h3qHdlgZMCIXRm9EF+A9MNicdLm+FVbpx
Bgrf9M4wsHU0YMn1vKjp7GNNA7IRM3msANWqYR+khlTMNoV/PJ7hHJq1C82jI1O2aVMGbrqHXCEg
ltPIqdulnCYWGxeiR/9R0Bck6FoFsSyRH7dZ4nSg/UYqvWcVSS5JygTUw8m0GY5IwhuCF/VZacpW
TyA1QooT8mCWTvZ//dCKZUCK8xZxrewMCFFH4RNX+SG4ShVzcYUMJBcsTuwTtVH/fJTU7qgOtevO
a02lsq7n+0f21FZDvfgUHGbPkMhIQQ2k1X3Ker6PH09nXlBfYALv+kZdkGwrzugHy9RqmHc3G5h3
sOwm9ZFnwH121VU5c/5I5jVvd1VxbOapdXhZFaZVHi72fiLYcxuX1rOtY3bFz7gTo4UxdmMbudRS
+zn3lSVDYcWvF/3RXBVjakgw5OPdAQ9s4kCaEapmPzGtJhoYrkN9FgGOcHpvCaVx3XBOjrgKkzff
Dh/sROpewLlh7T0Pns4k+5VUB3wubHcbDNqtiNYGDLk076CC4O5MOO9Q9+vIi3xk428lWBMGZydT
U8bvwLtPjMruBrirEBhyDo8xlXjwcSp4JR0wMMLOwLlEp4KaMIogbaYp17Ix4On/FO9taMVPCfeu
KjOdmmXU89J89j11nA2W1fOYLf8fEd32ga+mCxnLidLLhp5QzmokfckkDJtrrK0Ycg2q2Ln5VN85
GG7GrHOtRabFI+CMgHhKNS7gFTyDWgI30sn3X4q3VCrZhCZC5q0x9qdg1wfHuNHG6+PsuBHUPqq9
EBH3jmK36VJjW8Y9GwAEO9Q+I128FAATJaMLOd3MJ7/xj33MW8xoUR7xJaL8jyewRJxF9Lg701Eq
Ai6+zVVSy9DxRIeUuSd20U8Np1HW9xB7JznPv33VHhyWWgzNNZd39Wghp03x0Dc7zZjbyf6qTDCS
6B/JOBJgy5ySd7D2ANrVpbXpCLNF/QIlCddinNfxIPdmiUtuiiGP9830onXF1TXmywcqDGT9hwuP
NebHT0JgofhRZCL+RPj568XGM/qWPSAjQzyKKjIGgvA7IxSy0TP6pbXExjbHDha02zWBxIu1u+hW
7KBUr5ynzp8m0b3gDcjqaDwOg3lzhTQK3akrTyV5JAcukr7avvlkZELWGzcANWvmOuPcFodiEU0R
hqGMrTgloawWg7h1yVGyqCWS1kGTyeeYOvgIxkq6cJU3MR6+v6XKv0xSJSEn7RqT1exgRsW/2b4M
6Bh9C3kgKo8PSAPh3FYN/bWLUjYZUmvUoMJfgj1WTkADMmYm84ozZbJjpdlKQlrkOKL6ax2kbIIB
KIA3qZDozVcJQLSc6IlMVWGN2/hdfyBFRTLX17y4BPx02ITRyBfuzckuub/WG9EtnpV8wHWO22v7
BPleSqLW4GGO+uNcCrys7xRdZxzpZ+4eytjIDOWYSpXCc596xs+bmPDHA2RNmUXBcwrr3badNCgO
NKnRQzYxE4vAWo6b9g5L5cYkvxJp6G2CnAfJGSinvLxg/si9a0ztlQeisDP3MJJA5bWWKGwKHQmY
zfLkaoX3+3ydLgv8jOBwLXgjXatu08/5rTv1rXYbNJkbWONZm0uXzfordn8pg9Hw5YdL/nn5k+xk
7m1r1EhwTn+nV79DSOJZ+uz+tvXsld/QrI1RGDKkaCRXRYXVe7EEQUMBbP+Q7C4JKtQiyQixNpGm
sA1ZtMWGytxN1w64xrS0TSgisk9ZXmN1iHkWCS8DvUX0XWmEfeR5MmYXp2+nk5cNPXJmQlwm1LK0
4Q6ZLpUUz+BzYeZ3wNe16HMIRkTYqL14RG35Y6pnzUVixrcuxmmjNfZblw2u/82Wv44wl0P0g2jA
hqzIKIORpLIkvmLUsmSYILewhINpevgS+xIbvVJOTdX0XqsJNy/GONQXy/XVoxoE+PC4mzRfDtbR
YdutsmcRmFhwdlYbHa2vqNBhf0zx9L1+MVuBvwFojQ0ZuGgVE3Z4N5XRbOVTqnn3MPHbWek6SKBq
9t+G3gNziVye6VzuAF1aCVvK/piNn5UkVI9ROySrJPcAbQiMNXkZu21uNND0KP0NoXcGO81w1Yd6
hFCUFJB8C1HPwJb2obca4ic2fUDe1DtRKkSH3ePkxP0f21uVz/NXDSHKn9T3kppnpoRzc9BWyo6K
2siLge9sYz8wG2VvTGI0jM8Q4svUKaIXGtZhqCFbOHJbxtEf5cP1gS30shebw71kW8WhMQL7kWOZ
QC1GfZ+k8xuPfmZCSgsy3eW2Mw6XFSBfpA3/1nte3RR6EvTFl5LkIWBwKkAT1+9YkYF0q+isQFKo
UfKBC0rdvzdBD1BLkIAv7jANAf9mpRY3tYiYhFMRQR8PIkX7BLKwuFX6onP6Gv+RrjxzT4513Ueg
fz9r7f4V6LFzL1KHKs/0Zq2QcSRP7U5v1eUIEXFVN6F8SRZEMghsg28+OrLYh7gzdDrqCBydK7Jy
M3W3XheLIbzD+LSagoM0usoxpnNiM1+irsRI5zvtulJh/l1NrpfLB2O/UH2uBmDWjMRR/n4QsEgJ
OHya2tqrFdstDqG9IU9aZZxR4YoaaMTlLBORGtkzfykbilr3A42haqQbSvaAy2I1mCxsZCQ/ZRBw
S0hXHL34KyEQYnBliaoEByC/2Jsk8bClmAb3T3bPvM6lYmSGFCEvDB0ljdbWuQfMaerUfUCVA/Gb
3FvzbDxHKJd7e9ROb+MaJDXqO68dRIMELrVTZDjdQozYg/HuJTr8/ITEleqToY5hsAk5My4S3RQe
60Vpz2Jg+6zx5IDqVyCVlDcsn/mAf3EN8wNIfPMl5PFCg0aGc2Vti3SdxrCrthT0/oyXhN/EVP/Q
1FPuq6GIXij74+iTAbXCd2ufaBuFEOWWh+T2B/alAa2JPbdCWoP/wxFKBssXJJdj8auxmdRzzK11
nRF2I42ZD5OmfDyNkyZlQYQCjLmJ9uC7mZCZj8MnSxaBrDxBziUqrdAvi9crX6yB2GtcbgKfsWCH
rJ/iUhfYuBI8RZx7mdeqOdOxD0GcIgKvFisvZrVT/Wxmwv4fnRE0h3BpEbNDMlQTBY6HKn6JCuUv
QPsAJ2Inc8khPhkLfOQV7BdIrv0qfMo8u1VFsBP2s7dhuiztr0EQZFvnfloQEkXmf0dm1DKPaq+W
N7sD/qlu8d9+g2Kj6B53ncNrADv4tLjHzx4eOn3oerXGCbKxzS5FhJ5elNio/O0ikShGVi/eg6Dq
0s7vFzWtQrDi9pb5Q+A0zzrcemQY8Wg+MI39Y6OzPx4BHEkftXLDGUDfIzkWq4+H0kbrXGVZ5X09
W2UUskHprYccxG6a3L+/uH005GshoHwXVxWNjrOKq/oGtPpyinIZkCVhL1thCloRCrQIV8afEqxI
Ox/yojWYqOMpf4xXXsI3xHWsuJFvmB+VAnvoeQJR/27++uPzTplfgri4rjqPIMKpAHDTdMVEdzAj
52pAB8g1yAPlrOsBgScUQVr0QuZuc8ycNNZUpf2ZX8MNW2FTEraYCD+6YfJusWwN3d8QYS0KEE82
23gTT+Tud2YWWIQcb+EjR9LbHLJsC4wUjVuHTzfDsvPjcGvzquJpanjVtM5bvRjHTu2V4llVM5VI
/e/KVL8GxNph6tuEerDBpj/UOPrZaluJyLrSFKpkDtJi5siSX/8CEocSLsz1TpCqmJ1hPMbxnaaU
gZ/avBcGMoMGRPn7gzRbR20aKWVm0HabPJu2RpOT1uAtc5ftw+XCdIBgcYFYSWqXWtNf01sUTvE9
0BOiHtoT9298qQwhGuqf514kjqVHxBaFvs4FcVqxQG3h9t+E2mN1gyc46esPELYR3gMXXCA9Od0E
66icTMUt1TDWt9ecqIBXNEUfolJWWClEAugR2Yjcp1rWvCvSCTRK8MZTVS/+whIjj+IRwJnTouVE
PYng+9nRX4NnUhTve0Vut+EqFQvR2C6oxagnrORcENKcz+sY+4urPg5acRza4fbuUcR3R5Y72gEA
9BYhY6/dPPNKSGu1+zenrvREx3VLpZJUsfW7wrQrgBuLCT1LZTvGr/1PA8o16rTbcT/ia6clumAi
yOj4XXugFh/2AQHzjJtSP0ljCOWydWa9KeuqU8B8cMOcfnpgQUYsnPT/3DpgUcSR2BDRSKoSHVaF
JEzjYpO9Sa3p+ZzACSNmfEBsDXQ7mgeC5c9QLbQ8D0nF28LgQLDRMVRkC6FRvFMycX9kOfp/Fh3z
4j0afHLSSM3hDtG+bRA94Nu06fFsl0U084d8kgjvXtpeDvvjEMOKITB6vDXzpX1Ogo6zfU+KszTs
k8wzlSbRHjt4PwYNGrFBz2ItqMroCX1uYIfW8JN/qtKEplgWPtcaFcjOYUncw3x6Xi9j4kcRXUu5
TDlctf05I1VuxRSWKIVPkmMiKs+z2uUvxWR3fJrDsGVgdXPEPGyzyJ66DiZ6mK33Y7+digPSIsGX
qvV4aOgZcP3oByIgcFelO2FLXfwXjs6ZIYTNOeNajYayavR6GWeI/0aXbqsv2ZtHNIdME0iSyspv
vbAEqR1gz/QhVHUiMmzq7/eLlfjtf2vpD98r9TzBvfpr8ATybmRIoSqHUaDp2VLYR5XqQq34yM1r
hTfDsbhETZP8SIwu1lIBoJcqR90CVqMAh22EVIKtujNm74HWnO9/vT4MNaflLtXPXceo+/cgh2s9
Y08Dhhqpek1E50tBPqSeVTL2HyyHTtFvZLEIzGU10xMXZI16x2w4gcWUcc/+B59KWgkT/747QPW5
PQfq4ITBvFi0DI/Jnk9s9BVvIYipvXMLITSDoB2dI39LjYwLUBJvwj1BU8KMgi1cnaO/tfucfDFv
FIi9Y2IEYw8hdhnGGKTFZCwZwFqd6kvcRRGLJsRZiw6p3FLUoPBzPLoUUqwmYIF/+sHAtVMW0bqW
7Q7teB2o+lk1UsDrcjh22QwuiV8GRtlSsYQrB8b321kY/sAVAHbrzU53j18RUodTxwY1Ph7Gb/EP
OuYI8zN05y8n0CdKEhn+oU5kKdJfXLSFH1RwGj7kv88xhTwGuTRrT4Q1h6FHnZdybgJh75wsx5AI
QK6tJ31JdghHk/biivS17Fzq57toBDyk1NMm1GkZOUm1D6m6Z44Xsvcbo0E5KjWTFQuBakWInRnd
JXkrKwxrs2kYkwMtQ5pbfD5BucyAcZD11ttUKWjMYPuo/XmiIHHgosKUHKubamrU54u784vQl5iI
7IFFXSKk1WJARX4W5eezPjVlGTawqnNf4RJw9vvXmFRVtLgbJ1/tEk1d1bXv5HB3EADtNwXn8nqf
2W0LSWmBvnzFtPLuXu5iwnEJdlLfVEO5SuuUBrw7zFZ6m31xR8uSuojAbqQichZyimiowxGFnrAL
BvKx49c9URUhi4WDFnQvzsGkDBjwRpXQfPxnbyeOzGAS0fA7DKg0OJpXPvPfE28A5lkDernUupP1
KQThrRVp4wai0kHRwaP+6vViHSSUxRWS5DEUoJShHTav4A5z3UWKjqkqimrx6Fz86T1UYWG7B5TG
gEZ/EPyykFdtOyeKY6+CXki40T5QbsYK3Y7R64wkxZhbi7QpTFVXWEk8jZWCj9BTpdH/u0Z5x1Fk
hqCKRqA4xdLKxjIZwpu6d3YKNPcMpxjYSLa/X5XvTEW0ZheALNbs3GP3gttlo3oS8wn9WCAQJTG9
gXxyLolBe4wUI2K204M9rcFWkuiFU+uptoKX23mHBJVm5PZgdz+tBEGcWQMHEvwYlVtZVGsNzZ1w
npzhwnh0S2FibfDVNZFcdYusAxMBBZEq6Ro19YV8FQtJJuknrSAspcVBbR5/eGvzXQ60RTTKUoo0
kK61DfoMjjUq9dRLgNfzWEc62VGsX1AnOOb8fienOTZSkhbNbdUR1rjDOaxiafAifqGrme1E+wNI
kYLXZPckt0Xg9RSuI7eYkIkRrRQp4cqSWJ3iFalYUDIM7vWIu6ZikummUEQ76sJTDA0Pgjo+dR+t
+smTL3KGDeeZIHlvKn6lEGT8l2r5z3OFDeH0pMfm5LBFXZGlZv8RSvKy6e7jLanABw3pXFLfIawj
M9+tZhaFyhIZEdfsQhX8C7bPValcEIY6C3EMtw/CUdzaeRoLQa3nSyLmOsmDF1kgR/CgXbpmY+eo
E4EqGIFuE0MGmc2qdpBJYeYK/+K2dqqZnUp6ONJzzwFqcNnDCAtWJ3zhcr8MCfvkULt7qvb80Dpt
inGT1LBkWjR1GqkJ06GCxW/zZUxOCLYNIBoyS62PPAZc2icMzuCXJ/rwqOBisCptqxUi1r0QYcht
taiBR/4D1irzTn7FANYyvI6EW//IM1vmEXvEDtrGwF++nJLCPjGvyHxIYQ79acRElAv5HyMq1H7A
CgYH1czUOn83lXUQ4w89H7nAXrWml+A8Wrt757nPMyDL/R4sigOAD7O4UZy3Hm/aqp6W6ErZPAN0
Jsth/9dxTwPSOwwGS1anYR5iD2SZM0YH1kGkEqir2nmQrhdjclqiNqN9Ha+vG5N2Bo1Sosp78Lgi
KxR19c9vkQ4amW+VeYWfEz7MtrNpF3YQpfNdWcRQ5yrqlQ63n14ODaPsLK5MJhWGzHGLd+A5Pa43
ohDcUYBNkff5ZtvhsKCrDh/qV+UwoU/N+EZPEE6ghdL9UsHVTeSfm10lcnG6XfF4apMFyyF5Kndx
w7KkqOXNwnekQsct2bsnF9RN4/EcJzyHVtqskBRRiG07svM/OMDU3ocVgTSuEQU/OWM+zzYKpAcO
hMBUAthimiKo+hD1F877SANiW76xps7xf93xS711XYKl7STkNNFF0RhbFImmTtb5qVeeQuFlD9Gt
ex8XS291PxvdYowUfF9vVOla6brYlGrwmSDWhgr4FHBpjmOoLEhWgEF2fspUQDOycIyH3FR0/wNT
nO5Rs4n9s7bT3HGeT9mOHldbNt2i3m+WEFhIfJXjqlSXA0jbhWaTU6cYfEy9FwlmQQn4WjxwTfr1
ORJYxOKOffgp6Jx0IZhsR/7t6mK35Eks4eDJg4QbLlHeQlA6L2Ou3nHEr1be9KXhfognvWPiZhMC
5Rb4i4Ogd7oX5Cg0wd0wb8kNWOYLmMYf+x/6MMr4gAkVt5kv2ENxuzupRApwsj0Ft8TrvU8ZBuGR
ViU30r++v0I4G/sJmWHZ7Jk6VcYMCRAA7yx9c85Vq+LAgv8LD5iH/aHi2w1frk5XBo2Kadwlsy+C
iHC7pWW2Kfou7SeYNfIS9+GDfCyalI6/ruoeobyQ5CCOMDhrMWGrNVrQvYedUI0zsgCxESZOS31t
3LYd65JgTBuw2AJKJCRUiwRHCb0ZbP/8kxihQrg1Ih+sLpaUv1eTPlQcgum8pv0q2kKhsXH5Ifig
6xDW5tUcddtcRs3sGPknD2AjYcMLZV4bnjcjfZ+20hQttUL3Ey+sCrGOC98fDCsMHIYXPWDpbBW1
XjmshZ2g7Opi/9oFBAvDlIjf0PcqRa3BzPQhFmasboBGpV/Vu1Yxnuh5IFtVrvlmT2cEfzOkHYbM
hEx5uhzgcEgRFK/rf4mcdJXSBhcoycQbkEQ4Bh2TSXY1bO3b7nnlfe3upXs8je0QxTfgTSIpHclD
nWuJ1HWnqhh8Bp/8VkUwDeUJzTlTEjLI3SVyk8KoWEzwlaO+PDG98GS+z1Zq0Ok7SQ8tGdAjfQII
BEeC+pleHJZ/GICyHUQSdRbzdNI93d2u5qjS1IrXOfEckcsoiTdXHLci5Jo37qLyrMFvl8ffAd5+
B8hEfOSSxtLzIytKzncEHmQfhTm1NIUbFc7pz9dGINc6U/0dHY01NkeSA5/t3PWyhF+8uZpEMrFx
CfSv6uHt85NUjXnnWjXPLT3TJWwnODFF4Pe0hSJjVb+ADBt7yDMAXcJHVhLlWLBzpMdTrw5xCvGF
1hzuCTH+CFr79m/7mvwQv+IgVKxUnQwJUT9TsLHorwZHcVCvfdDx/2QGhuE/MdYg7ppYt+IGiSIC
QP6HfRzBs/47CWi0pvhmgIeiikuWSCkiyrg0wsy1gCIibLILEXZnmIdUA6CJV1AYluwrYWqTVggS
9qhRGZ0frjwubhnQYCUTG5Wuxvh+hEGpRjFVFRXJO/0h1YGcsYwgz82EuMgxnlTI3oy0wFP7IvLJ
W5fV7hQ2qn9z2YNyncqS0agOqNS3VCLnP3FSomFrVUSlw8J1qhFcRjN/YLu7byNbFmq2ff6uY3nT
eTPnhVAcl/oK8L4mpaPQ11sOoksPAjq6zKtZZ0qiaJg+D9KEwb7qddgypv9hLwk9dqB5qI6oo1ml
a1OwCACdDvm7OKwD52m/kgGNSDVDCQ43EJN8o666oGRDL6E7biQjEudtfd2m8ow01962UED83sfF
c3sf3V248Hv/YRs11PAawYKum9o3pMJKQv086lgoegIcIGflP0Yi3OHtvzfb7AzOOO7kaH4ES74R
Bow+Yew20mx99xuc9hmU71OWS6YdFcuT+ROw4ZamD7ljbUG6YQhDxt4JaSiznkuPEndmE7HMw858
T04oiN++CWsL6+8VL2nWPb1EnoJzrxZ5vrTs5o+09Dm+S1H/SH23s+/uOwOCacPbkJoI4qMDT4op
cD+99jSwi953IYTGjGTsBEyW8GYqtykzeFx20jw9E4iVGfx21RLRJcRNg731fgeK9MBqKU0btWji
GTwGyj3YiDZDwxHOcSfAeVExI1gebAaIYAlFIJeAn0xTdRgGHygcJbasAabmIFPgcxhbf8fffu1N
Ynblo8wOORrCZ91W7dbqo5Q07isrEsOip8jdznYDjPipmHLP3g/0+8XnTJHj5stxDHde1GsCinLz
C0gpHpbSslzahkkvhI23QIWwvQjhPYzFFw7lU5KDW07Va5AVvE+4OJY8JPrVPxD2qpbrdBuF1PJK
vEthvDKyzrS3jw4tqikx19qK7AsCTSnayRDKHY0kBpCs7GHNX5hNXKM/Wj4J0rY/pMKJMniQXQJ1
g+ILEVmD6bDvAGxV1ZIMPJsC/bITlvxTt0xP1BdBZBrF4/Z+zdAZsOQMWX2UH7HomYmmuuC3RrFR
BZTQq1gR8lmx1HyXYT3dTS/PgYCwdwsrCEAjviHeRCDqjY0O9aUCMsmtiZY/BPKFd+H6nrDebqiA
UZhT8i9bk03yalZZJK8hI+YwQEvp/uK40skwZt32ko+LEyi7jNR204a06MEXTa17lVFwsY8E3ZEN
eamEZRY/mqBTTyKcFSHBMdpAEvSYMu0IuseV0jeRofOux/fe1lORDohAdnssIvMx0b4qGH5qmDV0
UyDxUxl9k2ryqLRYY//335h2gm1NriU0rTnEl/Q5xyryb1VL3g9sGP+vFwJ/KrIgSuDO6ae6+uqo
QV0N+fQobCugPQXRC3Y7TsUdvgJsuY/QUk39yXp84D8wS2/gslxFfZb62aOR56MeiTTFGjzLa6H9
1aMB2v/5xcqXi/3ToZfbreINoEq1GV5Kn4o2OFd5U28VuAj345+kpFL+5BiptR7aUKYppd6Q+GtB
CJvJtsLzpE07OSj8Pbc01Gn0/yxeZYuttnIvZRVNkoG2+QtQvCJuRyH2+2P2eL1MDc5ra1peWQwe
CUizqCAj/sUn7Gm7RQLqTtBQ39GwqO9U3HINdkqWUh5QPjNkm059lx6iTPDFEnPbaeDWmTtD1f3A
qCg3Kk2JZ7p1/Rk2dDsFOd55eDAIYRS3FVuY6keHI8J/u1xCaSXnds2H5dHNtRxW/1hHYIAy+DC5
8HocVlzE7GDS9u5bBmXWk/RmwcRbMe/5ZwDTFpqKwaXq8Qx8Atx1glGC8x/g2Eh5CNQyAqNqi1pf
dan7IjHLe7wtvw0agrkwnGv+q4CaPrv5A2wDmQNMRvLLLsjGJV8m/SKwKgsIBNGPAaJe2b8vvHjP
uQgueUE8QvGBIwnSeQjUqvv3OFVOyqEMRsyB4M/cUNEZUawsnW01VFBlDYKoQ+vQ+MFYz7XhUfM2
JVtDZfEfT8YfiNAcNFrrUbnSXw/FtWoM7MuLhDbYoA5lfgsZBTdVW06MxNX2BIUMTuREqrySmnJm
5axnK3b4OzrpZkqEfg7MOZNgJzHiRiB6cnpEbs1g+S5/qg6VSxAzHJhWkl6RpdPbfbKRq9pwyX+H
04z5u3dkReOMvE9gVCuSO0xX+kPqbEfkfhG7K8dfyb3SYswHTC9M8uDwvcDUUrSG7SgolK7OB+Xu
0jgKRs781HI6Nh4MAUkwAWJmIU95mbVb1OgvK9H3dZGzXvzI7amY2jRt7J53cjTHpwY7cMEGcZmP
GoOT6oLDb4rKKwvDIAgF6ous6qKg658wrrDpwOlZELLQtqW7WWljqDtv5/URyKCeGS4usPIYLT7j
ceOMk6lF+FzHSNJgJU4HtemeAhkeiSO3uxnanyRYMWn2+OuLJP9Em5swyRzFDBbwB+HCvQWgtd4A
fvfw2qfenuuG2pw9WbxvJ9b8j6o2urDTMVUgIGIlB6TQm1XOgTDxZA4HyC8CPuVR+KmmAHJTHKrE
N3Tezew8Q/JaTGCCzcxh5yOndbOZtN5sXXDHxVT2/b8773Ui1fJHL+C5x4yXqFkZMAxrexJ3pYtt
Ic0POAUVuPclcVvbypy2ostUGNjxdkMljtq9f/WiJ35/50HnrRpvss+qgRMfbxJo0TJwG4N4qySe
imOUU4umxDWzgwINlShiqeLZGOgzHFuuJo7qRZSCrLdr7dcfY5MO/2WwFKYf98l/doonPKq11/hD
jJvr53dAE14Lcmw1sLhdHPnPASwQq60i0u7ickRtL1LtLjo5XpJyVW5pHMnkWGrUkG2HVRxm9a5w
XNrRX5LpfeCgAOE2MUx3w504pqH3NU3gScZIQJprkHdogzFCrkPUzDcPU4/yS8gXO9Rf6+LZcaMj
Y34XEVAuEG0n4Y9wjGy5xUINg1kPak68QJ3fXgviwVr1c4kl7qFtUTc8sOXt/JcHJP4oZQZ+N891
xTlMSBGdSrEgqdTJZ1kiM7nmdrotLQI0Bs1Y+TximifBu7QOVdrS8OwNcld4KbbnmYRieFtxb/4N
o88Wlx8LQvKbvoSw118rwcEMBYBFfB1v8253UGND43qVgQDRsBHAvXr09De4Lv2zoxUPxHbNAo2J
t9Iq988LYHODYuHH0ai+mpw3sH6maiG7oISPr/Boa0k/Y/SuEEy9hoGAomSWeMZJX2JtPWtOM5XI
WrOyLbywmNHsJK+iaF+/ykPl/FDKZyaEaaicmVCO2ooOWOEHnN7WoK8itM4JHJ1sHwtarHf04dW0
w39jOaj0ptGxTS4IFlmsJFpeMpiPDFGhI4TLMDQ6KkxG2UJGYtooIiiM02ur0S982gAbv+qgW2Sb
XBdr3wxu8Pjn13XcpOSamXW+DSY2kP7rEuZpFq+USJ9S/m/Wdle7o6m+VBlABGo0HNl1IYr/8bYp
Pgr5z2GZe3fmwzv2ZMGKzsCLQ7NXnIWAhxT56+/xz4gEx7cxeqlFXNDjkpftUjAHBfd6IireaHeu
d1zu+DdlDAbkGkZOBZomb16kvCrvBp5pDIq+HW/yCCDklHKEBxL3/Ko6FkG3yx9O/5zF/azdRG8R
Ks8JoHMENaEyFHmDYl2Y7h9uM+gO8tw0nCdGp2vUevDF9q83Isf4ZNx1cx2sKERw07mupP4DgPfM
v4L2saQ1B34AhshYe64w6GGRGbBWShjTM+6JHp2vcerlCM0r1PNFJvslb4UMTBRjHbNAz70PGv09
4TXsDpooUmInjdKsp3BQNxamCoNIDGunJiTXAmo7jbrBg5hpufGLwBLThCX5HzasCnSk85dw2ed/
u66BUMQU1heCzggIwgx5EZAOGKlDZhLoLQ+wBJhQ89jlr/BP9q9b+m3/s6p9oGan1Dey7vISMdP4
0bNWaRzz0zVASRmTDTKb3k/9BQpGsSlhiAUVJgrvo1H8uQk0DEr5GE6pGndB/Erhc+HFaTRLKKbj
9J0uAOMbSRkrLQaxegbxb6xcHdPAGlIFmjXWPzltPmlrJOVMsrL+JSSfecQSK/+FbwzdIzt+XkLk
jvV4UNT1qDytAjZRn0uEsWHzkWoIjBIKau5+cqWl/5HBW7seXubtLSJvOxKtZRQj6ymBLPv/YisN
+69nZ8vKk82SwEicAmKLQHggg4Wrt10qcZ1QcKQHV3VegNbPnXVZQrRhlckoDZM2PyTgR56V1ex8
rU9DPArzp4IRWGNWUMQV3ihfRjNCiq+sVGp3V5LqgDj7IFWZb6hijo0D6ABnGepPz3W34adeh7H4
CeTLQdk/6VOtGW1iuavT/HrAOG2yaQl1gUpEzk9JTT3bLuHVM9qt0nTMp/8lWhZBpVA+sl86JC/y
ajb+8MLbAA5xoMLAw+HGxfMLN/2nmh6p+o6+vCes/uu4LtnGy9CAMwcpXkxGqeWyva7zyzeRNXTQ
3nSTOecfsJCNjFLzX0OK35aW/ckvt5lDnxPuR+e5pYMD8psOEbmn8fq8hihXLjNEOeANpewiAVqP
82OVYV0Qd5kln9Dwzwpw6CCePZxtpsvdnJ3YtO25WXNW4OA8MACRpxkMjzUJjshR/mZ3cEY98PoS
PIx7P2GKDKW6bDUd7/aA65/FMUQgsBCGaDsSBfWZ+JwATJj/h3d+Pb1vBQbtP/eq257ibg94MIpp
OMz8tP/6lyyzZR2EnYwDQh4D+R8BuAAmDNGeFdPiKwKQoVwWrZC2jWuIm9YtDoDAkkHe/MQkMybp
laiUyA4oOvyFiJqgOvrDVb/mC9364oIiBogK6o27H7aPLFhO1al5n5XRU38nn7D2Qvwjy+RIqm8e
Xp58f2TmSiezU1LFpKZtkI66l8HB1E9l9sjeQHNudVvhLWM+WZIG/p+RL/X+lKMdTZO39uzpLCm0
AzpVOKh5NEeqBLCVVmvKBgYURDmLXh8rDt70vOnU1qpN/5/XbgbhK6gJJaPeaxxkhAXxMhR85p/q
/WavsbMzp7V+0YMw0i5DaatW43LkAYoOJ/cXasy6Masnye8ffsXZ25fGTg5hp7+QP+Ociu6lBHxo
6rwi104iS2m5lkesE86SmjgDDQAxotj5WOX0wGCsLfsal5jJmbatvQBDy3D3NxqKjP1bfmSi3eUi
QqNgLVytJWE2oMSUUI99C1sMrtlMOGsXldm19mpcobygQMy/OWddF+8BQ4+vcdINkkt604oARbi1
RpO3WO+rBovHuUBRmfNYXF/AQSCEl0kuIoTv7SXpqDGfbmdBo9knmhaoz0kr717Lk+ox8ycRu1VC
VS+gwc/vSwy8qj2t0PMME08hGbuspV+6UfTQrcnDOldhe+HRujfZ2i94vyPqFvILqeYnpLYxWtIr
SEJEGLi8TCOtk+gRlKW0bL8+Egx9Hmyd48prWKtcAh/K8QzqT+5KvZ18Fidh8TllPngVdICsgMvT
WyQcysSyg+xQ6a2f6BV0v/sWDLQiVfygkqxaL/eandwJbvLfxqGiAYmiVgMVCrx/i88UauAnJ4tT
XXsoTg0I+E8HwGQOIB6njA2ftOzodo1giTjmrDcDVsU/YNimZCO33AgoqQM6JB0zHUhsr3QDYYl3
RxX4Fi6Ek2mKKmc1TNHEyQCapQcDkBtJiSR3SqEVAUQuxR7kSz9NJ2Zifb+W2j7TmzSmv0kvYvao
LPdHKrh0vxdj8r1u4fbY1TpKRqJtcxcw+VbdtLwd4DqW00KbPFJ743rdPuDlHMG+d0FSr9HiJz5j
6/zDole/f0mCDpWcH8XoWyM7N/4cJqEa9i71GB9eJfxsrGyNjwfrWOk2GvIQSesxppieFqLhv4Rz
B7jJINbmXvfkTO3nVUAFlIyNTJPLWUu4nH8JeNve6TUFyK7ZT8X5tSTeSp3Lvk8Igfb1CXuvvm28
F9QGcSeXjqS/brU6PQmzBtGsLWn2JQsfzYH8c8iKCAyLS9NmWwbbQCOrRbDp3BvaUioM5JxRx3FN
Npk5ebqq1rcxih7pIuRAnpCcO48F0rD+xOimXICLeCMTinsEcpYaUuMNVN1ytx5ZnUIKClYKuG4e
iBoy+IIFfw6pulwOPA+5dAjHJwtyCSA5HymY/oF/71KCy8GggkMeAODJrgy4jOpXt9pR0B5aJXDc
4odMmkN9v/89EEa9AV7tNtewXFhlEn2XG6E/q/qnGz+zuJbtgfS3yuc7MSOsdcF13tifookc1ts3
oFDq1xpjgnMk2D+1HZVUlM1bv4Cfk7mtcjoOV8nYKZEzK/aHakpp1eflZZ+f9SD1kFdoAe0bCCin
DKXd6GJiOa4Ep4ZWldvSIPezGnAQAfxZHDIiUCfFw7wuWNsrDm15+KyRuGDb4b/AXOBFUxkJVMmi
eHZ/sVRd9nwoHGMmCrzKVDCMoSnkUDmppkcJxsG+EYY0Xpse9dwMBWS0orf+HbKP6fvUcAFJpWls
sWcewuriyEiIybOV8SM2aTbv25X4HxbaRvAqK+SxthTrbmXy1rD7+EQlBKMMY9vKvyc7sgsol3ei
8JN+ZcJ3YgKz7stQXLCYC3hdwuKf4qImehlPMZ+iiORmT3JxyCCVCr3mkbwOLRBNxckCFHyOpX3r
T4jQkO6lhMesnLlLL+g8YoO/gQhGiEqm52Zovkr79iRFREZ30ZcLhmFvVR3GisNtAUTa6y8rJELg
apICVutjVUXpiQCqLCKY3fimkAP+2gd+sr+KIJ3IDYDFHVz03iTi+Ux7bSjk15uYaXChJwbdRmVO
mg2ACNL4hDfBqjc+wpfQnQM1wYCkRAKgCpgOCC2HxxLIZfT0gX1Sx/GzzkokyrGRHP9tHBEbVKYg
e3JLEQn6q0PCOlbf+IfQQ+qAkAnYTaBUXo+u5QJyqSZNRkbznglEUnbpz60tlCqKp1vA5ia16F53
6SvY4altYvekSo7Ak+jGrdHUUgB6Vd7eqkzB0zRTtvwMSDUHRQ50wTuDZ9N6F4CRWKOmErxin1ts
GiF5S2zF8d4ywUTVgXmIa0jr7ZP5P0l0ERE5MTuVo2ID2Qbm5Okwi1IrKSZrQbosTYS6MII7lfFG
ei/fWYm398/4HjIuYehd3YX0QcS3+0D0yLjKIXJiO5Yw+lH7pffg/xm6CV3BwDOzrpAqB1iYvENo
A1hA3UY6AE/HtQUdjmr8vOzODsOfHKPEuaSQpoNDAP+pN0czeQ5LqIMlDmFPfR6H70NsgA0KnE+P
jMrL+S06/O7CGtAsPOyxt13YzC1Yulsx+BeLSXqJyi7hfTMx3qLZIV3wf/2dFBcUrO3Fn74tci5W
ab3w9lGb2Giljc2auWrKZvjQSg1q2ZZtNXImQMiNfJlTomvdKduN/DYwsvh86t4kYvVRYWp3QIy8
oCqyXufflMk1nmPsn34nYlO7hYhr4i293HwVD3fEy82vQYAFYc2lDW5eZnhg2b41ChYQyeH1Ch30
oDafZM4oqlGN9P1/3vc5zJfDyfV+vaYs6xqoyZCmlW1KnQQfqTefuLM0ATvfoIwB/czjVwbRvk7s
vbT47mOIsI8aXpChHt7B6SUn3iCTuQ0qIQEi4x+n4TTICktRVRsxub0mHhGGPuR2Doqt5kltpZx+
ZyBSoiaFSNvitgV3laHjepdoNi7VsyjnXEd1znYwedmBjyNSnkI3xKoMaDPIBozEfCecdeENWAds
sTfJey6L+Kz0s7f0ZeEIEXF6ekWzTwvb1rghQUpiPolGenACw5JQyWeFLMe+caBjruw1Kei5ADeI
lG/cyyVpTCij9EtYMZVSTKvLELJ3TB0uZA6d6jnsPuVaeyAOE1qVbTRoEnCMKnTr4L0KDXkaj/3J
49EHmwu9qddpquDDlCzGFt4jdIvJ7k8Fgc1Ccw8CmfSByjEPG+sRf9SVNW8u37eN5bL8iOFCLzqX
ZRxr9FGLzwMqz6xHtSfqX2ovuzR9p7LytEcsBIROhc/U3MDYtmZznkn7f3MekcqP5Pxoy202Ax7l
UT5Ju6l6OAmyuhH3aXZksO4OYgkEMgOcHpXzxHJkDqC7mPg9OQvSTlu+I95Cnq1uKzt6ObrEWu6W
Ksl0EPoqwfE8slCqToXdUp3ZE1/p98rDQxV1d/ap6+OqTuwYaGmly/wRHbY1p3Bmvw7Gb3bVXJGu
3/+2d0bpn1Gd11HjqpAEcs7yX+uhdH8tNKnX553whWVNwrzbnETT7ZsYRJAN0IJoYvmJJ2+XYZjy
fDFiXpqPdZWIxS2kATxPagY6yP4TpItqmO7TLKUuwMW742wdOQCXOFIeW5Ny6j78NJEZ4dctAIga
8Q2V6vluiCCW7qAq4AoBUwTt6QHwAvDSo/HZxtj64uRkKBC0WSkPySfwUyEKBJeXrlg3fMyU8uWm
QIN0Z5WPE+2liRXmV9wZJPhP4XsravJ7u0YE324iuzXwwW+bMTxRY1zzwAO0MFyk6BTql2pwgskl
VLwx7LXAu2GlAjSJJsCGKGCjO6yDiBrBVUlZZELmdAZUDSDODhDkN47Tz3hTtY4r9KhbFYvKAmpD
vjDuonDBBO+DGQB3dWQcQGT6FoEcXxfji5r+yW1u7ZOWhNwNEUDHn09IgwIrNCugn3jrzCcjI5Ze
4ueEvAKbQ0qI5aRMI2XDmy937cxxs6aF6wenzlPe/8NIatRLNwUZpEHpKXyxAFQSHYVtmkNc9Wqq
fgFwL8we0Gv98+nZ86DDwta75Lps7joD7F9uP1Q3YREuwlocjaHaZWAhB83hkQ6vB7KP4IRAtqVK
IYwCWjEVFBDM52UvH1A+3CiYspB/hLL5FiVU25bj+sKac7mWaXYFFqvmjpEniLIqYhCackHt644j
dnOdmUbfOQVFNkBDEHdT4cTpBBEhG8D6YZeZABOiaJpfEkxzqEnWXPpmd0Sas3729Ol/iPralDgf
059Se4hi4ROhWpE3Y6SbKdTdV2piygY/kYlIoY4pJc4to0oiv5pHIMUfKV2mYUirUVfOzcsRzflC
OyiLcMrHrHSkvww2mPxRc7V7Phuih7tPv8BXd9BGdOO4Ws2QxxMzHlvPaEXzcf0EoTS7I0jufo+D
ClCiekedXK83t2mB2aFiMpuiC73Ayr4FlIUDq66P8UFRSNKcVcZ8dUoTLIuvCbCqPTPzL5XdrZte
3Lgnw47ey61xjdU7doQKMC3hkMsndCWoL5mYME17ys2Yw+v2MK4P9GE10l1hqqOPepKegIB1pHc4
0mQTGYktfVdvq5U1oIzWPoRYVA1EAyLiaWeq6SCuA2V64UBqeej0j5dHoSBYn6tuX4/HzPLd7ljC
kfAg0jq3vzlq4lkYTlgxLdt86hCoBz4cl6DgwhZBye09ZdHNy/qpNQdAod7TwIoIrY7xWpk/x20E
5laidnivFVdQcKI8dAjKDfxR075Fli1di1lC4XeO/70Evpj31AGbTnDyMq4a8LbwEMrBiYOV08Ai
1WVjiynZPaoz9G525j4nYzJRunIUToqft0HsO+vdLjKfY1bn8Q3rjq1a3nmJhmsgq+zZFeLhciV6
3S/KhvmFbxMOW/bkL0rEHXGlqz/46sTm2d0zOsHTH6i9wmm/PDq1utLBUXnl4KxN5ZvwotjJjvNx
IT6lp3EtLaD9dOztujboX/g9zLxiNg5uBT2QRx3h0QGwekFtVs3sWK6LFw/p1YpHgEAWhcGoGaEC
uhLLNUgZx/aZbxTD2i9GC+DlLuR2BAZUM/jcwkY1NId2/pNHeR8U+DJM7Zvkgkq2GBPXz8kmQdrj
/rd/n7Ha1hF9m/u/jdRD+2ecc+x0HdX7Z1Rqjh2VCeo+c1tN5/ZwKIm691EFVkCHaGvfSgA76l8j
BJ+/iWKVogiu+sI3CHhBDhwvYWY2fLnlNke+0ZVLrd8X9slvO8nxlRHMWyhq8FzjVDvgmvkmo7jS
GzVK2D6bTJWF5kaq83W/7CoJvtPiDkEQHHmh9vTcfhsE65OSw2uzkaVMEVG+DK4KkdNHi4wUJ3jJ
VAkYu9Kq0+57im5dx6o6VJjMeSVHokrwx32h1kPEgOU2iHqRvADU4RlBd0JbUAp1O//5BT8SkDyu
iCdthbMdlvA1Vax9WMRdchkQbvO8/WmMTYLFYV7MA6dB2aa6myKnTf+98RDVnJioE5aMHzTPvP5A
MPno1AiTgpspnUV+bXN1HhSSA8o0GcJdOHVFcCV/9y+MWAq0LxStxQ0TRiAcy0PpPt9qfkVEGJnF
b/k+zVTYpSVXiqShFBREb5agDzKpm2rgZBQBEfSW9Bm3P/rnxOvtbqGJVERqbnPkua6kMbITm1tV
ZcdUHVOJLmMj7ZTbtAIZGRFpH/Yn4WlZwHv8EfToUFN2DjDaBFZFeSbyFEgpR6Io0zrKzeLkwX1E
NG0m+pJmGSMoa5+7xltQy4vpYCkZj1ykGNyjppX/ZiEbcbFpwS7C5DE4bnnKJ9EUhq1axSzWIDTE
xelKd7n2q/K1FdUgTTkJy5HXaecucH8rJX3tUshwoP/22izZzNvDHxBSWm5VCvm66/73N7XKF1Tb
loi1Jmd4/6EYAXrUqEZzoNTkK2l8yrScOZiwYxsqpwIgWmUEeAaDdyeAwDK2I+D08/RlnULDQO8V
FYnxtydftcMYzQH+iqf5VxziyRyLJcKRF0h3XNl9KbZc+5/lPf4ianwduxjaPl0NgO9sScTitJGg
Phq6pT/CoadKPcoRYMJImpuuSHVBwP1oYszAAa9bNNcmhad/DqHYrSwsc3/uPdnGQwbDIrzWBqLw
5W1t6x7OYYggH4xHy2G9P3ZqvURoql6CEOMm2BnLWfegTwU5JLoJaoYLC8TPOwWEOtYpbZmOcxmU
6njuWmP5nGPlZwQCjqLIzQeIzoCPnmAcmPkDCfGKKHbGiY+Ix6WlrMngD3iJf2Sy+mzZCBc/9sTF
WeZPf2xblRCDoAyY/pIoovqa6sJpizhUQE2JMrVlErxSS/ZrbyTgPJsCgtZQzuUeroHekJSDvRlb
6CZ28f0IS3OaafUAX1aO+ogMKGA+hNZ2/qP1t6PD7tkR/wuDLj9DoYHNVoS5AI4kj2Ad0DOy+E1r
WKJEqiOyVxkaJLJqQU4J4NorUQdEBMilvmfOj8TyNJvmMnFMNxWwEe5vlLnZT6S/9P+eN/3sTC78
MZ59m+55ZfelfrPSOitYudk+DKaxpHKDZKP7DCmFKvrgrD/3SgwAAMmVhYZ4zRo43e+szV6k4RsM
WGzV2bILVPWHESf2KXgeR20l60TcLz8MqZVo7X4MJfASwTENLFgUkRW7Ygj+w+qY1wrTgmSvPesx
vr3eL9sklm0e++FjvQfbSPztjrDJ9VzUfMA/R4mgbsMSBnWRVB8uf4a+o58JRJN8bwF5n0o9Qhh7
iBdasI+4H++jLkzE19JiTJibgUQ7gPujnnc0gjMu9ksQLBNYXkL97JThHQ7vFMfzsRhlnN4nBn84
mkgjj8JyMHWhFql9B+HT+rqgKUvDyMKoW/vYrrpiIXqVP4gEb03wii1yCxxOPI8jnE6V1raezgQ5
Rh3IuETm/DqPQwup5HU8Ow/6g6acFY8Dmftu8er7PaswAdCzW57A6fedZ9JwMNz6b9yF9aU2gbXC
lTOM76La4lxcm4p/ABBlCGHQiE/EbGeGXEwZE25DuWJyBC7CBNkgXeBF2REBy0R2oE4gL6+AWQCy
gVLO9oMcUjItp7fSgp/RrDZWV57JikAEbzvl0qSVHy+1qGjXXLauGPuUCNMTy046F/F1wHoifJCl
IRi1l+MOTSenhJ08vuu94L8z0EKKv0843MWpAw1XIF3UlUmeioafrFCiDnZtGIBg7Vn1xfBhCmfm
wSXloTGWUG/fAj/2rhtY58FEMtCIeQ5FoNEy7h89P70WPfV6tN/8iItoPo+feQcVZFcJDE2EDg0r
x+UAXvjFzPk1EDQX5ed+p5N/CXBOgw9ybA1ed0B4kfW04pChJ6k1Pjxt9THrbfC1U3WVhI3vewTT
eLszvowBTaiot1z0yC8WUaKs1s2SvRnUHZ5rBdhIHSumZoBSw0gw+ajFBUsTFl3Hf404AYjvP6Gh
KgjCIO5QXqUIeIblIDlBbj/IthdpkU3tWUcnfnIs3lHMp4bUiSvQ+U8rw2Rhk02dvEQx35GVXmKe
hJU1Nhz99rZP/OyX3uo2+pPh+vDma/MhzLKrX+f+yz8SA2VDrb2yGkQnKTYEHZFaab6WOpoAQPjD
mNH2zbcsppJ+xi8pOZWqL195Yh7A1/snqiM0tuoUY9ix7kf3YzW7c5Z6QAe9aW30rzCW+KayF6vd
nqANP4UgVVObzbtrThpzcmhhp7ybPdNRCnjKgwMP6XsaN4Bx9Q3UhJM9F9BEtUWphZfhQXZI7hcO
OD2s0GJIUicLqt0BruKWQvgfHIhBnauNT5xXId+Iuq7gHQ+vg2xVkeg40/M+4FwB311vQBmLhMiO
U9XWkxXnbyUAb77w/vCVt/Mrf1rW5t1ekmMfFrcSDl3Gxos05kdcUoJ3oenYVj8OhL/WmVmmi5gF
BoadyPhB5pRcZtHhCl11VfHCF5+FjX4aQwiqgPoNWIx40jE9VvVhSCAbTRHsKKEY5k3XGSQjjgg4
nDEFEMsVmz7KlsrqKf1AdViJJmmkKzdUQL7aL/JiIUMwAxDGrzjerMQqEQEO7+6cwDfz0QOqtHMQ
SR+mqypb4YitAlxC9jNBMloUcsiGIpRAPsNyJxnj/ROHwMkkpZ7V9xjv9TcYCVSw8a1MZ19bMnQo
HchLMswk9Z8oOPKxYXvoKWIlI2wiXXXmmYaGux5gfJHqNOynXA/3YY6kYOCDda76/ERnPYAxj6w1
g98F7iFVzexHXRH9q9O1cJCfm12tHAe6dle9zPZ8Iu90E08uQxRKVQxo31QZwShvLQUvtnqiTG7a
xDquE6GitZiS5nln+orztqNVR66CeZWBreSh8xf0ei1bthhjqHLmEICV+zSIxxgS5uyZymQs66av
TbskkKycDe8tslhoB+rlzabXdg65hb9FpyzoJexP2cBBqfpkqHxizWJ2svFmIIQewD2bkFUCMX2C
BNQ9jQqTIE1KRSraNLO/6lZMTkF4zmi8AeYVppw6yG4YdGvpI+EzaqwgL7WstvvNfFp+jGCLPSYW
Vka/1C+bS0eQZjZcOhVF2kEnoINcAY7nJDS1eqcCH8faGPmmYy8pcqIi7vQcdVNpxL7IhUgGGWxY
WvqlvH0twW3M1/uEETLcCjnRpGhpz/g9BLnDGOiVXd3D1epvC0/chYkJE78KII1EYGs7O41XZlWu
KCv8UZC9DRa0bxYLs6LMLW5Y5CE2vKQ094biBuyHAp6pp1E//P0W0TmAtowf1PnX7wkrN3Z89hss
DH+t5RfKFO1OHU5tpRxt6tEPyrowJ1CnIUmzIc0QZ6ZSrNoJMRVAAz/7XAbh2O4bLdvVyDWFJ8VE
skqU0Vxyh1l/pYr1+R935Ya2PT124FV8gPrymb996f9d0I8b3j0wRsq+cQ3iHd7j3p9zw7H8gZC6
KsgDz6hytSceMVrnh7jQKKkcAr63ky40yRKAYz6fsWS3i1mFkpiSMOnL6Tj+9iCdoi/hCRc+0XBs
+bWYs0dHeF4l74nFJXq1uY4eIJhz2ZpTRI1jEfqXh74QNbWA0cnnQifFc0xQ3fz6pCpESmqpkz/M
GVyEiKRf8bYCnuoICwaGpaEvY5lz15XIuyVkG5GVye/4/QyD1vDgAHjYvJ35HxIyRIWneK0VqCrU
5I8AqrKfOAXBxq+by9lg+mEIyu37/rRz2NT8Ar2qWL1rP7ybW1EoD3FUbhCIqPbKoqFhACd/j7DD
l4/5oJIVBSISRa80B1iTTMgGEFrycsPcRY/fK9dk4rTQGnBiuRTKYy3Jfh5OJhkwcVFuQhDYRKSz
J9gSe806c62i1Yhn9szTPiGQu55ixjchJxXxTa6Co6L5/5MIS2CRJ133VXPW3aPV8rOySMiHtJgA
mdmlsUUegDVMoG3PJqNMWOVzLu2VlbNvzuMnqaCcR3LCQ2iVRYpNXkt+XdT3FrjPSfiAbN77mmX/
6a8dgKU3tJX2R8rFa9LcFATbSuj5PM4oD0DsxstCeGKY0GzqB71rhUTeaXPge+8Zk2TKTnYZTtXq
05jU7l05Gcaqpt5UPpNap/P+8RFEVFZBVHdHwujGFPCWvtKXYvhQVFF+JsVAu8xl88UM3B9IdYcb
A6BJkYIMosrN1PE9P45GEcwzVzRcnoTcH4NTqlcWwiEga/7EbjNHXU+0qGZQLQwj+XUs6/TzA9xr
hYPGrYqoKJZA819hCXWO21+F56EAJ3mVvir40KwhJcNebyXUJmP7K2hC1G5D+Ga70BliKYrFvK4P
fasOKhYKnPK7mDvsXSkfHoOOfsuLS97nMyvJzrJgoJZGo5ABfn0wyEFlW4TfaU7ABYhkvaeFTFIU
KRKxWX6DUPbLqfX2d5TjQjbOPLGcWPiRDqBlKb6DFVRsjHmikUD/jbFLeRrsktPMm2wZisvPskUd
/ZKQm8ZqyEojKnPskxgZI81mM8AgtJlhMyiIhqw+51Abthnos16jhhUoEERYG3j7NFZztQXEAtYT
K7LRMsuGqea/RBggcX5YJiuAK6QqmjWSc7Q0Q/GAKE9ByBWi8I0YWquvlUGV2o7duS/QbTIu/500
LK5wLoA5oTLPirUsM7hg6sT+DE9DE/lY+LEaCxnbu6xYB33zCZma/D5dD4mLfC/YQICHfg8tuhYT
e7XymXbG0HLm4YoAKGvg/+MwPjC6vVdPlVlB2z8X/DwEbCEOGTYSnWKJvYnTUduZms9wzzLqsEzd
EW9tl5FGMbgsYjTGcgBML9eMj1vD6I+UFKVrnifS0soAGuWL/kGvBDSnxHGcX+tD+s3HKRluksUm
lfBtI+cVbnvqmosctslIiVKXhIc7Ur1nwQXK/PnysppaMLM6wGacWdoD1G/mi85xTEaTqQsbDILA
dvpuJHUv9wwG3BBLRYaGp7tfVFcKnKDBgwS4X5WJ4NX83G7jXRFY5KMbEvyxWtpjb0ppEjUHrTvi
3ktLrmoXOmw/hSawpzZwFLajLyUE9rdw1kDiDXGYj1whT5oCOx85sESfY16HnDcpXzuRzuEF527e
Y4TiDDvIvGVWjhSTZ5F+AXkRo0d9ErtNatGbXprC+dYkBqJ1XiVOR2yywnp8BjS+eZr4bWZSoUR/
WAUDnlNFCq6K5KZ7x3gYhpxXCGeWJ/f43MNHh6glZFqe+Lxj7LOZFbFJMDcLaX/dVvzDmO8YSwv8
9/1HwtTgIMUewfyAzrDQrH981ZIrlCtiJ+xAJ0z0IkHO6ghPT+bI1D+2apQhu18ydcaUUKXX6ck4
5SSqcYzY9iUza5x95bj4S1oanMN99Zn02vBIt4wSlmm3DfF8VRoGoTdKpc9PpyPpdsAEjDdRDnty
PeyPbaYoiWcvFEqgWL+vsGj5cDWsu/2wexrHnO9649dfR05w5jMYkv4UDJG2MilPZgn8pDJMuPLh
+rdUbbE2RmA8g7MthDCKL08UYTM5ndWGCiFYGy2ZiYSaOk26gsl+aMve6om0ca2WPzo3ottIDh/i
mb3U6TUNUG6J6qiqkzKCy0CMWlJJ5MtWEi+r5uyCEFffPK2nptSz9QhOOXdF92uVwxYxPwNRB82k
T/y6bsh9KOc9thZnVjm1AsK5egKbTrjd+aqlZqdZKU277xEvj08xeMoptkM4JSqeIxq/9tUKgrRl
m1m43ocdKF50ifafhLFYf6RwMNrr2qjwFCuKGO9OS1b4R+PTGGDxdA41eOUFvICHyEIGDyvLl1lg
SlWS7rY64BgFbrd9OPhHfOgjG8Zfy7bVSvsphyuNFix5bMjqGczp+BWGLwFJgJJlxzwGFiaVhHke
DzM++FnQXLigPMWYakwFvSh00Y+crgr09CoQrhho5EOqD6zDq91/sr6uHdmBaaCPdRz/DZ6L+W65
YEgyamybQIg7HroZ+ee/7MZQyWaDs1XkZQ36j1Y3oKgNyWf90IzBp6TCBbOgR79o1Xzt5ivPp+l7
zL5WUYerJumozjRPQFdoNp8fIN4vDDWRDKqdSxAZsv3na4qAkn1VGcRwFIASD0gzQs9CZjsOej1G
I5yfhyVt7QRjWD8c2jKFATHk6qC+FHkPGHLgBQ1nchED0fEYsA4zHNGFllHnTDvhN/HGv85nLKTq
V19nlJz+/ruPj2hVrApllyXjeLkViBjLpmNlbeVv/8vQoBWeQp7akcf8KMIyLimhgMjhxp+Gj4lN
lDIYME1V2qTFzzNgVjphuc3fl01KoCy2WSRcSdAtTiqiUTroaks/uu4H5VpYpDx7OthlIHdQxirt
fVZdVYEP7j+QUYQv57EwSmYhQ1ruJIhouJeWxfwCxPolmeElNQBhVoDbUCseHxhTE1B+9fWmhc1t
DRc8YUoad8vQ29e9Qb9lcv83qi/1vju9+i9Na7OEH5uouWC/fddCt0V0g7Sr/aOFVMmiB/81VmxQ
wQdeVf8kRy+3QGTKpaeX419hXngo9fQMTfcbjlqXeMRmXg/k5Cois10Lc88IUAd/XV2eIzLsQ2+x
lXr7fyG+6xMDV5PAXJ6UOCvtb5e9XeSFBPSeMyHmTZ4xO590pe4iakotAHsFBCRxaLOsZKZ224gr
L+nBQe8HJ/bkLvF3ND/yFnJ0n5WUnzeWnemsWOqmiSjWphM9uZHXdWUw+jqSY/s/uYw7y48j4mdP
EEMp4MtSYQGqOh4UDn3KnrKJUw6ODj05/T1fztQzN8KrJydJJt3u7u7CJLm4bWP5SbXvWg3BJAM5
9JAS4Qc9BcIfxJPaGVWjw8C7axK/fXw8Tdru5sT5IdhQdmc4UsD4gCeLJ04d9HK3C6a0ofOp50GY
pBgWMcvXsSeetvEnV6/kNPvyiBhFku9B8OCECP+V2w+PauPnEPECzVckC39oAMsu4CWT9/ybz7kL
ozsgFFYjrLsk5tyRA46ARu3dzkhu4dS9eUT1fyxL016Y04XkJm7sD6C9UbUwKsjs6cjBB884xQBv
lawCwHSaXisUnfyyI80oNr6x+Gl/R5ZfWZIZnXYjtPwPA+sRZr1kTzRBHWCVqFuosMWQNO86SxB+
VbW/Phcx9pEY9uUcyw+hzLpruTq9JyjF99kSP3TrIciU09b++CnKtFsyfzABYcYC9AAwmagjlqI9
ttiMG/2VaDzQzLFZcjg/IP0s+c9wzk+P0t80aEjn6gposei82iJdsXeXSplbMk73Ay85I0mpg4Oj
6/QSvNHA5sb6CPYO5Bq06gM7am/wHUajBsTFUYob74xZOeos1Z6phsyrdRXaNM5Qf7U0+UK13FiO
PoCx3d71Asj35wZ158Jetud86V7j8Nulp1ISAcJDi1XfpMkby22CqNPU/a+7exhNcRVv7HtNW8Ra
6RZpmd4ezdpUNZCDjvk9eEaGWLHDZ49cwmSBT0hLm5xbBq1uJshRP88VlJ8Kx9KH2+q6AWPbm+5Q
6yCRcKRQD3Iu2ItIJnVbHNOAYtYBioUh7r7YFO3RxphT6lUZGpDLRrHOfrY/kOdZH6TGXGOtK0mj
Avp4p5MzVwQL8vptUIFpZeYA4UF9ADVM0/WH2Rxa6iTZC52qFLtbK4OdnSfwYm8+iXvzW4M2GnS8
DPrnjQr/PuAmuYnwYYTeOxc6CGhhf1R7k3QIUM3a/vtsushb9qIHMgGpec8ZyBrJEJp4IzWo9ZRo
tTnjeGOEopguMFy0SU/gIsAaRTeWOAb4zZPbIWcJTCEWtQBO9NODFqVgjAuRskDN57dnB//VrzM7
gjqYSfvQPnyRj9T8PK/J92F7RYLMt2g8sw5qaCT3H4FmtQl9xbBh3J/9hpurmGHtlxMa+Ign/VDK
oVEkUsB0Wouq5RFNWzy8tJfuu9fsapKh9tAL8Bb4I2HnLad8HF3ALYDJGvBBOvRNnr730mmDCxrf
btK7oO/hQY5a4Y+H4u0z8k4OeWyulmhPxwG8xcfywkneIXTlXmPz53LR7WKd/opwsXT6a0GQjoYr
nz111R/igmo+o0VChQ+szfLvMhjeTjymaq8lriM/Abdog4VL9MK4t8icTZ9pmQ6xt8bnZeU3HVq6
koWXPe/I9wafNePt82ZQe+70/XdrQX+CAtM5HzpnzLqoOHn1YasNj9T/lJpWP5QOZLaM5JQB4Otp
kaLtNMXAFaMA3RqnxITP+Gz0nLrf5RO/JkYC3BO5h9sOiodFQaJ2aT9JV2PTw03or4dID9qeZtrf
NQphZLPPD2lD9aRAAc4YwBA1EXN/6Jq2yR1C6PjoT/6A0dl9/0OPbM64ej1Y6VWr2ogNNZm1iPwe
e5+J6nSDE8MFbdWZ/vRlRVKVxw4iQsnMz2/5Er2LKdk5O/g20N5z5xng8R1y+L3E3Ni1lHZpsc7y
x6UjdauWfH6WXq536njoHbb9BNPyUQHWVq+DrHCO7G7qI1+Pc5jaSiXhq2T/q7ozFnQQou/wI1iJ
jfFDj+XYYyKxIFNxhJXxo3u+jCqPfaddCoVhOQqtJG1qF8iPVZfJbRMJBA1l/0ZlYRVd7u8hVSeS
iokdNAHm5QPmU6aMPooBEuNGFZKhjedlHNly5wkoVHN9VqQi647dxSiVcfEfRBhuPqh3DzI9TZpy
59Dp/qVXbEMFmdqmjWhGwh2na/Mqpl0gxSJaqAd1Wk0Vjg9a6Frov+LKaFDNCOKb+DEL5LkS+wZI
0wx3WjYhCnzYBKR0lO5dfkZ2/CgONo0An/z2U9G4v1KFwK2h8khZp4DDOhgE3rfL7zkXThBrHKcT
f5WigBRi1ar1BrVVLp5GE/tC3by/1tZNQLom6ooVStE4irccNBWZRfDatLAeb/0Gum/u5EiG+/eK
NbP6xw8V8wislBVyTDBIwZWXzv740P1tw/i1Rb07wnXcgiEvlxR0tUIB3Jb1e/ZvU0rcDUE5Y6eo
A14aBzPdS/ZhO7LEtTRreh2wjvNGaVL0AQUr5lNyRlOBbl0puQf4uQBkoHg6u5MXu7SJXUQASNJP
4zaXZokdUk4yM/Zcn1ZM6EXBLaLK7npolJ1N3fs7Hon1MrsXUDPtFceGyvX4mEt5lpppKeMowRtS
eofE9cCCCibKqPSU13szHayB7m9J418l4SONgz5C/2oSuFQI/KU8gX9o6s4J1yJ092tr6rrf6fns
J+3wEupTGo2xwwqUQfQFWTG84B/5yXKwGjvMgdxUpzxqOF99YdiFPLy0UBo8Tu67S75LI7RPJeyc
PAkiLEJHtS2fSW279xaSHw64zSLSuZZPnpM/L3Gwos9IZxIdjnRrCaUXVdl8UUC9OAYdJpXyQyWV
lGhNTrH3yxL9CrbXlaI13Jg2cXn+3KdSVql8GIMIgi9ADAz1Rvhsg7y+bTW3Bnz0xoPBEZTVZGi3
vJc0FgLutKJHVH4aDocH5vhsFm6NEbgmnOAV/QeSdbb8dhRKtkls3+mbm9Oz9cnwgYa7D5NVuDtW
5M0U16H2GhnO5vmgkxbpcEN0FmXLuzP4NhIKNtLPm92WzrJoSWcjFmomUlHekSMWYiEXzAK8akeV
+KhJroBNrrg7qWH3WU3WPRRXvm77MQIjZ3TdYhiwsAP4WZVLH7+0aV5yo37G77Gd8+PhrAOu+jEA
WI7FtTJTXHRQDPlntoap7p8Um691BmNXzu0y2kQ3orkHWc9d3lOLjtGaZFFFrDWK2I0tbBs7n7Zd
sxaVwj/O9reXmCmpgt57Q6ztEUNnTMSnXQQvJGwkaljokY1lRHID7A/jfbxPKMlLDBq7RV9V54MA
WGEoszIbIOKAUXvPISl9u0umELJnYyTqxrSS5xdNuP/p9m4Yv7AhZtqK+EZ443hO9k2Oh+GNAhWY
qXmCon4DchpQuinU9G9WciJhq4rhzwqJFMOVScf3TZZ3KFhErccj24eclCgLCnaJ6oT/Rj27ho8A
woigL7BHaBc8/Z5KfrwuMD1mQlFj8ttj4W6NDcrtzoFb/IC3fKMa5adO0mXsNkXBMQSHb4GWGDwH
SoYTJORD6/eOIR1fj92znkwnD12qQ5bUuPh3MGWkcBtAaYese4Sn0dd4pPrwQBuRJ359LbUMWeyw
6q/EbhzsbYu0JBxgvHLSJUkD8SqSo0KhTsUxoE/Tgadfg47ZCHcHJssb1/jpNu1+jb0eXfA7RJkz
PUGEE6gCycsE7kSsYvAIGb5HtGB5AE+UhV/f4sfqp5JUPYizoy9N0+vWW5su+E37GJZRoyuu/qLL
5v83DWvGcHg+B9+YerROK562gG5XfUmP8gvFWJnvIPGKEDEOUSVdE1uwOvxdwHzT6sT7FMZ6/Afz
Ns171YpOfTI+d4PJwb/pBXs/M5QZjGtrn8mpxT9KyW/5uLH2dGsM9jc6E1pTnJqSLf+7yqqru+IR
XDp9RhDgHLP6un1H16Zhkm6/UKgsCSaLfCUVM8KnCkuz3uTgtm7due12oUzxJB8NdggVEJMlFEOI
mhb4tMBajGdeJan+NLaWChLvbKVlzQyVukSLXkoAY5xVLE/B2AKPIwDxnS/satGy/i14ilabwHLg
X99qW2EAgfUG6YQn5aHZy2mgCUV7rbfZMwcQAvSr5/oICsa8tNA6O0A6ySwDYU3rv1GW2tgE25ki
dOvFooAfbAJQxCQChM0v2zizgp+IK2sOCW4bwWeZn9aYlG2TPbPovZ0vFUSs654wdppx+sR/EDEL
qnwupEinACX5Qk/pGjo+hLVeyP5yYwr7vJ3C+6UuAy8esf7THFwRT5XH9GmoCRu2wP1dqRZc4kQA
eVs4flJKdHlLVG6UqMyzeqEckpu4RPEpV8sMx1DldA8EOnWkFrIZirWRVFIasutFlfUTBZUVnaio
Bt2pgeUKfOOZSd8oAOwBfUh5scUvs+4keL3CmWESg8ukVLBUQLgFVqaKuUx5kjnB6hkRPmODx+Fn
hF3YlGU1hnJ7GwflrEDAMSsIE9JZ8NUeURYNLo6HjLpBR6R/b1VMmemDKSCJadVFba8of7yQRP6W
BOVtaowPg/oMYMuo4tGcF/l948xskT167TRlimQftfJl72bFqJORddUTAa6m5Yso++qzGB4eFyiK
iVqBGI6t8gLvf+F0+IVj5baCOKqqJJeF59G9vVGHWZ17p3uELIloHaWKYPE0I50tOiiftHnH+CCR
y51lfg07lm50k/oYySJfgd8h4dk4NRFMSyGoWE81tXTV6KPZg3TY2oIczUR4Bk2wHEnL9aju42I7
yVT+4pq6v1LQ5reYUOAP/W9EUpHUh0+Aj8EBxSKUV7ILebnz5j1J+2yOdxkBoRsngltExpmlGa86
gop7mJbVHYM8XsVE6mMzHx83Xm6o3dS2hvo0zHJOVFnkQOsY34h4sleEhQAUiq7x882ViU7aCt2c
ahwgKG6GFMQNbeEZsOBI2rplwPEVqx3084AFVME88u9+Y9i62uez/vF+LeVRnahhSYWZR+jyrIw/
ky9vhMvboy+W2iCGmoZC/PCBH+aCR2XJs/rmEZR8NelhZsgjAEDe2MWV2Cb3r3Z/0tCPKNFpgK64
Q+n8hB82Pr5Wvwciuwi6cmWcleEIq8uPlRJy40tnilgKwm4syktwJid9MaqwgRwikujpLsJ5zJZA
TDC8VwsYPLXvhn10ryYL+Rdp2oDPSOrVJq/Q6sVUg0ELZ5JKNVSCPr7xj0v5Fh1//5OqSdERekZQ
2JaMlFIDikuEi+A6U3PQACXpGIcb9RG6q0nmbB06Ob2Dq/ozEUfVYF9UiK93t/bnnFQfpObl2CY/
kAlOT/svLygqumAqsZvpg53w6OFwkLGG56MkIQb3oUlvKp6kT3oe5IRzqx2m6fnTtDTzDSckRM3q
nr53gRTEXecTkbG1LdhHTJdl+RzETRnKya2l8R8Q8otWqYA47ta/Xdpbd3IcwYzHHxRaMCVBHRNE
3L8cX88xsaPuhjjqJJ/jTM7DeW4d2LyvMFbd1nO+HqWVNTGl8yP2KtqJG4QWUPrIW0pugjZZt0iV
8g/wntDmCCN2Np7hcBu+wjQ/7A/wfOpLbdYt4i47gmH3G6SivzsjECL5IOPtgZHacxzMmAw9ikn8
jBRGkyWkQquTxt6i2Fe7y+AoSIo48AowCXcsesPyMi+guJYr9UCWtAWmJrC9n/fy4buwGv29n8Tr
qAfjmwA/mqu96zJ7zLNyCgsRF9ZDRrHavRNkV2ujsUTNGbTgnrhG+CwbD3W/eIOe5pujI3ZeGRT2
+cWzA4WSfdliJhxVQYmDN/ws9U9Il8zQhSOqhTfvWAXdBzgSEFg52IdtOmh+G5wepmdDZ1SH+NiJ
T9gbrsaOMbCPIjBQct/hRnuAvHR9FuVPCD8T+S+kdc2qBxyB+BRhxQi2N7zKq1GYc5+LcO/Eu/p5
27oXjKsK5SeXiwrcDvTavRX9OUmMxcarLMhlk8SbZgx3mLO8t4ix7b1lgSa2SxF4CHV6QqfdFTK5
/4JmA04kXcxr6uMN1BeAudyAhXh5uvHy6SxJp0fxJqJE1QHcl41CIIGfh9Sbh37LvpkkdJ4KuIQu
EMr6p032VHB8JYrLKehOXNc9KqOR+UCbgt9hdcRXby217WZxPhY4YR0/9y1Z4dezRDnxgV/X4Iw3
RaFf6QQF7r5YRWWWHAW3XuBk2LuDS8qvikKqQ9+dCI5++0AJ/zH9uXBs8VMgJPqz2aQVBONb0Od1
Rv5oYWt/wkSKwglEP6hMSmjq7Lc6rhpv3a21ahKHxeY/j6Iz5TZnAyc8SiSbbMZ6cYwAHNeGsCZr
Actq94c3ErhUfiyxQDanteHcBkPdTBXwdGrgLDFc+BZg2AMJxcJVNTDfnbGi4iMzW3qJ9xDKIek4
WQhauCJ8e/4f0Cf/ckWVJ1onLO3mbtrNxV6tx5r6lvrKTyejKdo/raim+Blv8405Qv6IxvcxIWqI
p+xh03J6d94hhTNbsCeOoQ/heL4W8ImuDfNQ8NVWv0rswDGU7B9j4Nny0K/EOudZfjfNPwe/S5Rr
GUqPGUdU91H+hpEydq4Xw297U3XS6bZkr0JAotoC3Z2HzdIFTNRi13rhIKxACbXPOjwC/rxpSY6J
ueNOrr0gRFsmcqDMWnSNsAx3LIS9tTLbWiwedhpVS02ugTFFFcVif7QeQnrCy/N6qMNpFTaru87P
AL4m4LNrE0HoiJDyqi3n9aZUawXx7cvmPSbG24rdZmM/NfQFGdvfDwEfaOqL9JLbF6TfSV2bu4Ry
ME2MNeR3al238IiKfltL5+P5/1EpfgPqzYESfxmLLH01K5Io9WqB4i/u3fAJt0fCuVrJ59zUhUOo
p9HOUdgTOHL8XEyrsUW1U6t6zcsZatKLImbuaG372axRFO6MiKIGGxRB7zQNbLpdknWzBujF71ue
dh0Yg2TedGthmHnDZIcZCuwGssHDgDefnrauWwvrCCxgeIageXHWm7yzrO1G9pnAhLwQDpqU3Jf6
3v6UX1f7CMZjkkijcFL1YHSTpj2PoPePbg/mifHuh24ZTW6mxqdt9tQSmqwpmN8lxIVeD93tuWJl
5JGFBI5ldsUpt9rp2cRlkAd1b+ntHon5AdZNwamONJrQas+Y4gEI6kU8vc3VE8b4IO8m9Hwma9Gw
fSYXKUJRfPXRZIdRL0T3STOVnJmkhIf6UkrIlfFvxraOOYqdvMiBwmLu5K+wVXML+Hpf9s/vIvBb
xHd7W7qc+TL0/CJ/VTyFSzZuhtLAJCWlxdJOqrTHozsaPhJggw00JYGSD7urQ5KcOvnj2vp3MxVd
2p8bgJgZs4O9SOsM3iD88Yg1NmoRWiBp1VzL1VfuRR+JPESvuhc6IId/YwgF3gSwROJsE8x2F5/H
ZnEuqJpbcWMdJw163p2WUW+82bP6pabzWidYGEcMj/7/KJJiEgamRn+8cRMyImCyU6EtSob5WW5F
4xlj/JgLhxTwoygYYeerSDJl//vuNaoPYe+wE4TJLl3eCFSdeAw7Mz5W7UKC/CwdTP0rQrvkPNc2
JYsjL0ROx0aAkv24dtLAETihw6us6U/EMueT4glxnOut6q1yFXizuF9Q9kde48zYDnkw7kQkL1EP
9AlZO/Bzxtvyr07i7L/6k+j7llLjZ/b0c952TPU28ta/GYaz7SHssgZbQaq4mtaxWqgJKi5eK+vl
ZzUrOU6ecuia9m/WBMu51HIcM8LCOZJDXpnTV6REvOxAO4iI0tAdWV3xpzjHpLlzCCB+zBE1XFNL
xdnuStp0gEWYcw9GeXdXwuFT1bF4TDZQpt2SLbZiMgg8VjZrglps4N3K+Gx95z4jTBxYrBxdPkAJ
NN9VdPDXoeudt/cvMhbO99823O8Og2NB01f/acezMuoHRdLJql4P2Z8MXvURKtoEB/9MTQM/YAqf
NnoxZCLjZlnWahbxxmBzWQXFxO5xgOxOday0QgMQZyOmpxWiwWQOWBkQkWNTJbgcOiIiOtyXiGZ7
VLwWzPFJUCZUG2gYLLkHDzfZvZrLEYUe0m0oW3RFmI7dBEz/GPJpAXlRhgY1Vs3aIRKhhVCAoiB1
54ZLgxokmqBlpgJiB5F7dcIY2S10kpe5pgTM88Vef/F92rcpfpvZ5eAnzbTYeSWSAdmrso5xwdXi
YiD7L2otiwnk+I9tCAnztuMy9vtoqRQgGMrbCeRo3ez+VnAdZvjZl2CiYOYIeSETzKDWHP8XZpng
F1r18OvcszGO3rSQNw6yuPwnSGuXh6epH8UulMqjEy+3HUwFfhmeAVXXe7rdvli1X6sAuZzXZ42p
c5R5HcUFdKHOcDoao6dkJ8rmWYcladYWfomTg4BQKKLWXhy+EMbKutZ1V1PkdwW6DUqEdrFlj84N
nvbhJpIO3wdf2XJKXglq8VBEKWafaTlu7LBtzsbyd65rKkgfUlSQQ62ETqOxLir64B8k/Vh685Dm
t3ucle5MZlmcft1lSvPe6kkqg8xRD/avqhlrf/rbduPtMcxil+fDgIH93NGZbFhlotutyxTDO4tS
/J9/VmtbwHSl9I0rexndroLxCVuKLDvB1fOYUU9GczK3Lbscq82X3c4Zar+c5xii304DS/dTMPfi
ojOzwfgHTEd5Fj9wT9KypHzw++MYY3Ye9Wvc0OwbqpSJvdhmpnBaCsyQPbmlrFfuluAXSqFlQECj
pnCYYCLij/c9yXrIHy0YR8KDtAHcKTijILSHWeVwJXGDiiHNnUPo8bVN0nn/7rUVDEY4vDAc7tsA
beP9BmaPxDi21ZvO1AVIzW8hTXW5fmBL4uB2tz5gaG/endAC6yZcoud42X2ZsCAdWQbVgTY7OiJn
nI5PL7b0Z02dwglGQpbeuovi074g+6qfau4s5od8zjmJpPW00tS/kaKl87PwolFOenItqQqVVWEt
YzvvpANv3uIC1p01jbC+U2gRaSVS7dg97u1a73vsA34Q06QXsB38CryK0EohORCKsHuuV+lxz3Q8
43iOFpjH2NX6h2sp95fTdsS5Uh4mRqMWOhwyrTx3G0i2v97tvLuCNJBsQwDVUbsspH468F6mVVig
JUHXozvKMxBGW80Pi+YhEeoRZEGJsyCLKMOeBfUj6Ww8S7Ceqr8rU7/2cnREp3IZsFZV5J/7N0mS
tSAlDlOXvvMcb/vQ0Bfe1rVlY5ip1xbY3JTpO6g+Qmi0lhrF8oRBWL/j/hvw8E2ij+VTR0iHSEep
IYup9Fhbw/B35DXjZxJWWc7/E+Zk6fkMeqz4Pp1qb4dICjiJQeyAuMdn35LRn3sHcoA+z/0+PrZE
PiYB/MXT5vsUu4rGaVcj1r1ugkbpZiEJGEImYGwI/+3mgB5gZCOWG5Q4tAvIRe4d43wUD5bEYnfb
H29j7oEvtJ7z0pX9QQvwExzpb+Q9ztf5RD/81AqjnOZfav0LlYJ1lMhEZP2yzf0LNjygkUN1JYns
5qaH//dgwfzapP1AJ1YK5e88NLcsBmdLx1iklyTUb/zNoNjFCHIA/uT/ARVGH46W6xIwO9qsD2bS
9IPc4IuKkP2uWAIhgPEMqV9MQW0YEs5nf8ljOGZykrBl3iOaB+43SDa2u1QaWKn+2RfN0wSArFyA
gzxvEvGZNQ8jy+mvveemOZDT9oBzPPKsql5I2I0S5xXZaASe3xvcp3yLP+8Kpbi7Ija+MZPeuNYx
JRmvBaPoPd2bjozRc0ZOybFiXu4UQTW2xvlZhWNcRT8qrUFlQ1d6HEU00xmUYVCj4bA2bXceYkSd
/XR2PzISEMZJugj7DDPSK4tEx+RltKGUXVHQps1PgLW4gjPMjEfSBoJwDcCJdvdu8dUQ4fKoWPYA
xwKwgzxg6p7yb11vKBd3tYT1KZUyHw4oEdqV67TpIjQmkTC42g8ayt3R1F0U/XC7ycH4W9VRkRi6
weX/FYzT2ehjwx5fG4rkjAKM1F4f49UzWD6AHfab3dPnxlVVSnga/1iGLFTh/KUQOH4Qyx5Tn6bz
0CoK9qyv8io/oVCQxO1M29BQcNMLGy0/E8vXJH0wElZDw5/s3quQlYaYSEJV8gmUK4qfugPG+n8M
O8+FDf16M5gWoG0HdKDjAvAK+P6dWGwvQ6gGu/Grc8yjEw2AQVP382sIjedZ2Iq29A5pxz1sN/GY
gMuga6ED74hT1iBNuBhNDWjtZrcjYh0BzJoUt+o0Tn/cS9OR9XukQ+FdvsRPNuhIUyYMt0tqMtuR
JjiRJPDGYDDINcFTpnM7PAxTIY3za8edYY/0pSUN/AbsF6gPkF+/eF8v28pNEv8dnCe9wIBgyiR1
M0IbCc7aOzuSDU7LgfNdGT6OnH0uFANZYCJf2qToj+ngKGxMdk2nmx8oiaLSgsIpOCp7KKkuPIbu
6xp3zGYa3BQqdMX7m2/fMBqGbseXvWN8rYPJ92vyfGObGSQ08C9Y88UjwjKlG+0lwaxQov8X61/X
IszVBhcInnMTihR1xvEPXhuFnZCdyQhw2zCixl1D31cIlkwc367aM3iZ1/Vl0rw5YUbl90/duhH7
t95MkEr0dJfgUbLQbOAJwtR9coIzLUf38+0gRrJarFSq4diwjGYFLs0UEOfJDszbyNMGzqV9yMb9
craDwMGo2tqYs/hn3Fs2A46LsVC06hceTYfKyC2fBTbNaJmVitPQ6CeuNrTPXkkxdhNvSwvAiwpW
J+agXqHk7k7X43mEdxZgUkqti8TDVH5nu6kdeY8qJNYx40t7zaFE+zHPxBBeRX4Lc/8kauIzBTGl
hMpy/BAB6TZDyBwRNhsi9SWs+lOgyp1r+AduhppDEC1GnXIhMCigcKRel3BzwDab+rHGduc+Ee3g
uLSC3VdXt9B2M12WTtRuPRkMaCpnhpuzf9f28+CH0Imrk3o5c6OKKIcwCc6tmILZ9oxvCD+8dAS4
9EdGdFjnVE3kFgtLh5P/DybtK1dp6wuI3uPneEPNaXICUUIchZrmysRAXJFwaxye5idlNGzVlQ4K
7KK1W6bmMwL10o0IoafYjJgtYq7hkRqLgobgy80CtGEvHh9KH/OQ+kjPrBX9Pjg3/1YJYBjmcs4q
HaQYnp9TSy0ohmqbOWuvP9A5ULRkpaVF+L8sNm/1RxUdZ+AVgy7C+FfzJFB9GDy0C5en8gR6/VsE
wYi59qNdnCFMh+1wKgfYHUlS9GB0U2b4IPsvd6LDRUrjvbvh4+5HCEcQEwexFILjTz8HmqZYbbq6
XxUMFrzbxBls1QRZ0cP08XHnNFLopaASzT+ORQ03ZBkPbrsd1Ycmw2xDbX/iAz1vf0IzG6gA+tZz
/EdwxkbKYmHEX1RjaLgPw8pXQyfLDkv7dSm1xiXya+hcgEMwDcQ4q3eDNIgr5UshU8pgrY03kXPm
WM/x2tP1WQ6EwHyKkHC2zMtRbVO2ZYoDUQLsVJONnpnBuXnH9rCeevGc69+oFJzUDozWD4OJzqiZ
ub4ik5Kg5ZtNFdMXL4e61O5kbN1eZOGEsPalbpzIToGLsf4NN9BfTn2gGOoCQqQ+BEEYv/N285gp
4QGyk2GxJ34tbBGtULLUDLMpgwNTOldnQK3ilOG6yWItxEIFkxfNlkJSg2i1tyemxuZaRqpWlDzL
6N5shNiupG8IMj13M0EqRFUIPIc3fZkVaWZjybMJ4c+pSqbhN3TdGXR4Pfbuygmxwx8vym2uH7Yd
2BZyMC6clFoqwuLsIcvMwhKeOPTe9FlKl8jo7Xy9GCxCcuhVmjvgdOq+/44AM3mhjByjz0nRDI5C
xSHpQXvRi4LRUFZ6cNDVJSJBiA3qOGJb/k5jyue6VM0GQ1GrfVe46thUnY7v3IE1Q9ouJPyjW6Dk
XIGlRjIX9f3t+bWdw6xpPRPD6nGqt4ItM609+ewADyyObdFBorIL6o4NOz2+QkbFqVDzkjV40xRQ
975tOSzwCiZ+ZnOejoVK5hs/5EY6P41zMI1/DlR8bjzR99HKW0lQZcsgRFxObASRtKyzz7OFwdEF
YFcjmv848P+fnuTMnzzQYb1cljiGva6BTsNtVKdqxN77aeBjgtnPHX44KdrwuCDpgCxEpaE1Jw0X
MjxeZQYtS4pU00ZkFFJdU+IbIhGVQTmLM/6z/5W1DHJnB+FJDDD6JkehUKMVZF/lFd7BaBlrlOuZ
4GBbaIucBqd2BpebKXu25ylOcTgKsAjLI6S23/ldggAzxV85fFG/YVGTK9k6BCIukUIISv1PH3Vb
x1bmCbuvKXbfTen7sfxm/juLzMr84HYEk8k4S9WHxtS+9CNa9HcDtie6rZIIMa3yfcwLttB3DYFO
jMyg2ODvKK65AV9f6ThIiO0pE3ZsW1KZ8Nm+ejqWZRdtwmIfgDop4Dibt9ToJnQB/9sBLP04SpMU
uOTsU/3BU+CrkhvHb04qKxyZhgvsIaMzI34QusY7tcFn4AWJvwEKnFjythQiaP7NTiIb183g/Mkt
NvBnSrXTOTVwiKOLz6PfZdE5RegUmoVEAW1JFzCpFycvP2efWzF0kiHsss6/CNKr37JiCCDisV9x
u6XLfRMGCo4OxIx3Ypu4aFS9q13ZKD1AJCYgvjaTp8bsvkyS5FqewhZagv2eK/8G0KxD+wthy3K6
J9hSXL/Zl7DAfvNKjwXLWtsQ5StXVVjK0qgazfDIvCgmINikCPKEO1kzKIHqdqSYhP/KxOpmroaX
BRoa0RWUOuVzpMud8fLa16uD+uP5wE7GRNwqjZTYxoNkld3TW9fr6jHmyMoOea3m4Fde0pAlPZWA
OWKJ3mcRJT0ZaHC+J1sA2AMfcE07TDN2eHJQokf3UmglpMrsRgxtDfeCeQVjWjFGkAvtbIhrqZPj
NbPwS1Q3FVouHBo8J2ZSY/pY56ILqpnFAj7fDHLnPlTAJG0nbzgaWl/rP6+Xk0/ADn3Q5eIrl2kZ
GDV5YQRnEo6JC8GLMYgn0OVnIKvx0iW/+qqT8drXr4Z+L7AOEnI9b9Xv6omzcL4cbKaWegBZacNU
fMV5ejeGfSzYYfaTGu5WRI2FXc1xzOiP/DGx0HsFsn0yyrq8785yirlm25+TWe5h8Ywd4CLd8DTS
6brPAQDo9xUJerxVvoL2KpVDTSV+WPsfpPQN8GdOPhz1mgmSCHfwU9x211Oja9RTGIjDMXl0EAqX
lzRJYsdyN2aPhsSbiNHIfAgTswttkonBpZRozTAVFwAl6jw1gkvTJ6VIJyio/gvNoOAnOxu/gwu/
nXb9MUrU3NL9EktEzYuxt4OgpOrajIs4BYabie8dmRzrNHbg1WSLBPV3PlsUYk2x2W8F5F1tg8W2
KBv9OVuvoOdfpWea9Gb6jntvQjV8yzouAEereA/J0JfXr2wKU/jgKabf1ilnaetR3SRaoZtRvrqD
vTW8Wb3RJz1wd6XsvCtIG73LK7eHIexd3DbsP6J6jZ6P5K0QvfikMKRA2FLyYFXPU7gwCVwa8Mui
MAp+dMUsBi9wBcsC2lEL4nFkH+phOUCiqjRgJDw60fYWykkAmXwoRTQB2Lf+jOBkKOAuXri4bWt3
W42SEQRK7vxOKjv2n2iL4jx0tiXzG3BnyYLPFHSs8/v+Ge/KPJuv6X7Fe9t3rFSfzT0DMlQfp1Kl
k6v7m11qDt6XWIczIPx+DYKQdKrgK2MRfkRZI4xhFPCaXYiXF5N3nP7oF/AIanQsxHM782P5b2m/
6NgZHgpaJi4o/Q9P5ue+EmJUELDypxnrUgjqH7Xfv9+vnXj6b0rBp4mAujXMM5o/JUDa2Ipt4k9L
NoXWknnDWhKp5FCo1AcoFHVhMhWOxLYJFBoLr9bCf4nyvgCRCZExEal1DwAzboRVFHaBLyKkRaDd
5nkWqNx/9tlxjfLyDj2GM78w6MwuxARNFK9SACSb7viu1X20IPAqqtW9L+hTTC7bh54HCOi+epr9
CaEyC8imx/3Igq6H4EnEsYKUiCi/9eLyXIFv7laF/QeHRfhOCRP6GVNPNVZvZ5gy2DN4jmzyFgug
Hx2njSqXw5voynvGGVWsQVCFx6mUVst6LQQwZHU1iy9OImOE9DwrBHgxTW9OXxfUA6+VQNC7LtbK
l8eiRXOVKuS6FI1QulWxijw5A/GNTOUJVWh0lzYYvAKiDgfoaN76r2k52nWg/b6n+ae0i5Eh8pQB
24/QZctfkomQJ4V/mtVAmcKAUIRA6jUA3CeJVqPxesH6lWeFFl8USn4MDqy+PSMa6xEJiiJE0Xvu
Ub2n8eVB72PntmH+LgLt3BhsTI4hRjhPsemGzY81Jd2aNH/f0Tt+/zcVblf4Mwp81hMpIlmJNgIs
7F9HRbBqnHueodfbQLW7ARz8f1kwrXaHUDRtppth8S0Na4vnZcEkx2C5Ee9aLKW++POCp5KvDMzc
64/ew6XPyRv7QT6L0xjN+EQ6BsnoMPZrNPNaAE8o+C5b8m5+0Og/M8hmUcw9GVZQlRMo2dpdUEiR
R666IyoY9gZxmLKB1OGXdBP18CcdJMGVi4XBPlATIuTCn+o8VvyI77OjAqR1CJwQZyeB2gA8jZLo
kG0ExiD6tczES8txANZLpb4NsyDgIBVPTVB6VS2whuslW7odaQzlq85UZJ9MkSR5pLUliR4lLupH
tc/GWEFHgzi+s8CB3rXVvi1RYTWYtzAp4eaOW1JTKqcsnU+rG0spBhdhA6kL7NVn66ksOno70nUa
oKO5B4pEBx5bo4AW0XIPQaytCAK9bE4Z8Sv/X6q2d/faE+bpv9Mzpuc+EppFLRFToYoQK+y02XqA
JD+kjwPrxSyHeQhGfWmQoTYCPDHUNZi3iyEM2+CdNbJNB0aWI3BSF5n37CqBMw5Kiiwk3N2oA+PP
8CwnJHonaCuNyEnnrR0AGXWnk8WWdCyzbKtlC68BJcYcIgpBL54Q+/X5VRGBQDeurMp1poc7BjEi
mNezbEHsbw6AbfrQPU9QwkBXeR8C72/BiMyHrFWdrsDtYFFQQMvueDnve69mKULKPrRLPB97QkS1
cd5F8x5WMeTNYma6URjO1NgCLnXi7bF9wF87mjQ8mwW7YvePQzsHr4ecQSOadMMCagEboU70wLIk
sRNGGB9CM/TLPUKpRJQb2FboT03HLOmDT2NpHIOM+4EwwHOw8G0R7cVAY2LqfrNFrYBIxmWF7EJB
W/tj9prtnsmGZRafIyM/OoW6EgnCc5vF87qg8LBt8rne+VqFa4A31QnFlKdWqAqyoikbBlsr7Wx9
1TZkdL4SQPG2magCIeCEvhvPTO018HKBAMmKRVkHKFaERflHF5/XQImueP6tVJBfO6ZPcz8+xtmk
vSpiWdEMbtENe838SrYUG/Li3Fd0L6EUAybpYqxrisZRordLoVlmepg/QSTK5T9UP2pFl876Q88R
/zbgxP0ga4wMXDNaptB8XUeZfuZDHREd0Ytre+imkyHUXilWwdAcQbqXBjRscOBK+tHmVHpNST9m
Snol6shqmcyVJ0n8WCYp/FcKudn1CVwwTgfNiab3vyVXgA54b0+ZtnC/3XwpRy/KrZq2Ffo+7C5s
gMcNncNb1r3knSZ4pj/2jo0ArIZB4ulQmBUNoWDn0MlPJNIaL9vqp/GThsv5pXksxgrt1aXv82xr
bQf3JpzEEOGiTencUc6srMZIc2NuMt3QvGOyZT5Zo3c0U1P7vmeAe1e9pEDrA0K4plp5g//0haBH
GrbTyK9Aq4wOG/8ZmTgvYzMmjRXWru0xzi4xcxgqHmed0Aedl8t7zSIJlWpFTum5Anpg4I9mLrwv
WdTnrv2kaZUGySvVCaJIw4R8PS1p28UptbEIb7fPQhJ6aQw6xVAZHR1YEO9KJY2kJ0tvZmCVV6IG
6/ERwlH8tbpSro8GVK68/xXri7R8x3KQ3swdW9bcQvDQnTV/KvootnYOgUtsLPpIYwnwglvdGG0z
yARoX1mBG8T5T7/ZGc266ep0HxYBj+0sD97GK4jXssdD5aG67n56Mnb5wUskJaftSBd5DU3jE47I
AHaTTmrh9tW8fMABsCyrgUt98yRVFow00Ait1uS0Hxfx5adUW1GYDWF7WyEgUGvju/gmFEDmf2RS
2HEbygLyyvOionZvsI4e6EolEaxDOnpxXfSHruszWyAJudxBRG2A9GDbTdcJpyGFcjrjEProXcj8
YRuc9XBaE17eqyTifx1O3a26vkJiTeooLitnj5QtyAKKo1aEXzMB4Z4d/avuWTZZ1NvgCq6w8qKH
muWNDGlNsgD+vL0O/vkH1SNZdnP/xfJ5+82Yony4D9qVSpimDhNSUrZb95ESIJgwgSpnf0cc+z9n
yz7jTDosfRCziB3/jjouo425kkFSYF8n+kTjzRMhmT8kApVvFTd5eGGkl7RKAfVD19nPRXpl3yCk
gH1IS8YGJG3dm8icqWmlsWBd+zOWFpPNGAXvCTVIxDDVRBOnDakTvDY+UBDveeSiet/6N/zKhRJo
8HZ7RC/CZRag0K6vsE8FMudis/1FYrYN1cWeVFlSUJWpKPwW9LWhIXHHNmHPum5Sm4HIAmVurQ7k
yY+47Btp4aThKrIt5TsRnPwmbQiOCbcIbhqd3zPDlV9nNHqEEfIoWO3ANist6EcJYeMnbhfXNgLC
q8/6ZmH4Lk57DGGzz+dPYFZ479dV95gK5/UaK6QN/wEjI9YeGm0UmzMnZmFYAoGDYB8MGIjHlUbQ
z+RCHarfKWyEB+fL+pyUKJUE5jM1cC1WXR3NSqyNfj/ezOntYhChwGNWMuLH4c/GDOyqsVLvQcNE
49A1S4gZSBdFHeUdGKr1IyUJ6FpJEZarbN40NYpf4eFwxzU6dhEF+kgRmAIkomN0FK/RIOdOo29T
Zn86gO2JttjbiBOX/FuJr+3FF8DeITZYFfzRnVFuRKi1Ux8XSu1qab8p9H+w0IDn27iXPwB+0kvF
aTuqUBVbJyrdpq1S89/bFGz8sowgpNeFfrkc+GXUJaI+uKmIg103bAxoBZjvKe/w2HkM6E4yErFP
UtJugb+5KUlO/s0BfwwTShb9/ozFthkq90zFAUmL2GnXI/oSapgr1WpmFueSGXLraIja6ko6Dbyh
g7TM5ngGzIVWBeTrMl168zNGZ5F7++VZjHg3GloYFPBnR9yiSC3t4aZPvB+uo+14kEDEzOCL/A0E
h3dxs5cANls4SGzGnmGerpH1ttRWdOH5et1IVw9YCS/sFF3ND3SOVtWp3ULulCbqDyPeOs3UMgpu
w8/kT0XxeoU5H7Ermrav1qAys/s4dsDjn/UdWvgtZfsHRAhExPcphpyo6WL9jzgs4KRt7J63/nTv
A0tirot3A7ExSS694izraUU+enrwLuBg4nJSoTdadfSr+XqFSeVG9qmEJItD+mZ77IxlfOMkZWJK
b8+mRrB+TlU0liJcAYg5wEULRWg00G0vX24hw3MhwQo94VpwR/3f2w7hPCIW2nJfeqMV8IgAVYPk
qHSkIYtL7agRPhoO1q1a4yo4QmFfgQUXH/Is2GqteGWwCh8F51AIGprud7v5vneYqT1HwUIDRF3w
JRiytewwa44g60DtJhiossWmdZ/ogApw5mhRiwbswu3D96iP+lr/Cj54Z2zPdACjJD4P21a74ogV
VH/r29OQbMiUFe2Esks7JaN97IXKjQ0buENXp5uzvmZYhIyIi0I/4CGGH/oMCKkN5/t9FkPW/tIW
LJgTJPIpCxMDelQVLeX3JWWQwVoMjuRBgASrJI/K54c9VCfLEPfUIr+dQ8qXnjXshBwnJZ6ZUluZ
kWCz9ubC0IFTslwZyLbidW39a2oSYqbeuHTwPLsAMoW+hf+981o7EPARgwPl3cD2+eDpdGT7qLdm
giMjQAJx+kKtVEEreEgC7O1Bu+ZRgibFZmyGx122cach7eDjLNmELBr/td2O0lVe8oE3dd9BPHO1
NJ1DwkSj9SHqvDjfdzBFinKtKM2x0QeunzCvXgi9ypJ39d8+x000AkSphaxkjna6G26c+WOlFiwp
0Y2eb8G2B0CM0m4dFaSY1GySTJiS8A7bFUgraSf3dIkJDZTJe+fzgJ0Jh/jDpanTAVCP9J5I1PW0
ZUa3gkO44hjcPoBD+tcfnlkVA08V/wlTPg/Hao2nec7qGb2kvmLf+l8XjZaSi3Z5O6Mn9uJWCcaC
yCdX+ltwjp+LqLEJRP3/y2QUzMX/6ksRxljmWjZ8mrczXpssWRbyQrhbTz4oa+efRdRtf54M718d
tZxRjh3+2Ary3H3suHcIkYt5FXJ/m8iusfjKKfFWtv71VgAy80ScYhNh6JA/zVAMMio0p4Tf+qmg
JyEQ2kTh2o5c9pvXxm/E5GO68cbvodHj683HKC9/LH8OPFuNZm4h3ZnNi3Cwe4wirME2wlspaSMk
YTRmbkPEzGq2hQKIgUelQ6eW9AA6H9H8vnSra3lEVcL6KEf2EO+VrMBmDR/HRJ6z5n9OEyEC8a0Z
6+wXp9sBqW4acvgepNh9aSvc7X7bN91xuQ4lRq7uMgPDSo7WEdUMdF0EvSR+dmSzIw0G+ShswrE2
WNHrxnlZC4eSBY8oA4UTF+R4Fw3uCLfG8v3kRDo4Qa2+qI8g72KpFTK+jSwwvzq4y1KWStst2lLO
83fVy1qc9y3EWK/5tmUMWBu2c36q32P4UbRFvdoTf53E2N45JzT8DowIMdprTPNhM4wyzJ0XhA+I
6l0ZVhtNDLBFujk1P6ekWksFKWfDcwMoxfHxRaeSIdkG1LWaSoaDgMxh+ZeLZkJAX2wQOePS0vmx
we6KmdtW67KV8IqmkABogc7mLVEu4viWuuEyoN2sfeSTEsvzjqx60k537ICja0eDz2njSAsyg/gc
vp/nCi7FX+9tzUmwZ2/A/+eWETskFIy/8i3NBtGnORhFuynaUchh4U6gu6+IBG5TTOCigCBIyp8h
svPSNAu9Tg6FLsgaB3U+8ThDwwtjbdQVSMHwHPQV98menuq8neFj0gV7RzDf+uzVdIKVr38WrFX0
aoUdYYAnJUxrs2szLzVrW2wEWEH4XMm3OI6QLlpSGxIjwrwrxHaLYULsG0Vxk83qD/otoqh6UL04
2OKzMCaNEo3e2OcR9x1O1H8D772b8ZOBQgPKKDroam8QqpL+LzvF46/nn3LE1yOPUxxP4pYEyKQh
gxInOtUwILC9c/rtw8ntoH+7LQwRIvQoei5YV3yrCVERqB3XAqJ7o+c9cvnExt+ki9fhqmY7WlYR
HKfY6TB8c9A+6EWjj/gJuu7v1x2yi6I1X839SC1zoqVmUWV9wGSxR6C5LdSgIi1oWO9mzAr2BK4o
htDbSXQZodkbpQL54JblJwLC/XKg0c5uRZhRoFwy3cetGvFteiJYI4/pINs9WT+7SZntspDSXh28
5Q6CTela/S1sXFt7paR+ryUJWP9V5fyDZd7oVOHHqtRRrg1Gab/KFn9q4eqVBiIHX2+pGxZWsyrA
FQG8rufiUBvZr42gPTyVezBSzXdZ+EG/0wYSwC67hyvI679EodbQ08+wQwqOwD1i3R1XaUZqjzGn
hChXDx9+qpz/IJqPCXGiSzPMIlPi24Qn364CdLHH6aTvE8Nv6hKktgMP7ZTr6WQUnHLi4qtZHChy
p8+6GnqMUsXgAssiCHPPhADLtmAVZUQqiiqP1QjFuGVJAHDqb4ZhM04Q9EgRxmxd2Py/WBZmjvwv
SB+cCwpBWDJYMWAN1l68hS1Y1FVggqnMyUaa1ufoC+Ac1RWy11V0Yv87Dij1sSlGqzk8go+t2iwD
hld4+iZkqg+Jf0gTAnUEhM+k5Y747/eq2k3tnCjrjyfDlIVCZ2I+QOB8NUChbju0liammelyOzVU
kZlY2YENwE20TXjwwmjna6E6xJkmdqAi3RpVCPnFOEdxSJiGa0UFaRkozFDouUOOOBqT4+JvXPEi
584DIyM08qJb96NoFKa8rV9wWQeCGuJyq/Um98S/GA+QfDvs9R1iK369rAVaTCXkzMftx3+FafNb
WX3Dna7xb534CrY5wpSCj8pZEdLlO1diyw2/aC1ASDgGtFLOtgS81zG43AMs5bBB6UhBMav50hxr
f9s0G8PAIgIYT2NgmTIJKc4nJ83IPvrVa9djlp7v+26oXreJzgsxl4TT8JcwZWwbIHNkLATw1G6u
5wAji2tnxYyyGLmGpjyIeQmIRqZi5p/1DXg6/3ivJ6fUQ7AU+5D5l92MKZxtzFSibCFfqStoT41B
B5bUrj3gBlMqNGxU/cYKTEn5HN77qPedEoYNdIrlBVPi3HXYZChJyfz6WlP9FkC8AIlg5ZQIjYAD
ETl+xKA4A6SfWryOBJ9rA/kwmNqUi9gp13Sw9+A/zMa+ey59unzzXgjTd+4yCpvov/9D8915bUfq
y1W5tNh5yzjK8atQcA81OlA+L6G/6jW3VfKXeIoO6XMT4bUcu70tbpdiblH8LQ0P4Dasa8vLiK3h
G4wev0oSwVQdqMbtVEURXI8b8VQGTJisX25UH1AHOibLInxkhgarVBxDLZj7VkugdWysrO8Vxw3F
okmAyPXQuKZNk74upmt3+DuF0DRyry1xsg2u1+iJqWdceWlZTcaKITfHBHXRzm+1yd6l16LzPybV
7Mn9zXr4G8dqr3GKYqbgMFOmQ1guQGIM7p39x5FIiBmYH+F7aLorTBCFyCKiZnKvWPgab+EmD9ym
sH4C7z/z0Ad5QaAjeHqo80Fg/K4fViU23U7w46XfcxIAWJc56Wt3LkHihMpINhzMo4wUTESkXDKl
Nly5mhg6FCLMxhtjIj367HSOUA253sPJruAJlIo3CdcS7sK4k6HBJVvoC5Y5EAHa+oXgQZxwkpV7
WqI3FAqGvbK3P3yYZbBnt+RpPmC9tyw7BrhcyMGfVaZRqC6wAeuAunnq7gLHU8q/oLE6khQmqRHN
ZQXIRjMr1hl9eZec+jANZddtJheKjisnTT3VKeCLWosDsLgJz6ddfoRtkf4a79KZ9275+099EoTR
UHgLIqvyfvBgHlnxSCpc/uTqHA6FJJOKLgJMRd7kmmK1ZVjkwTd9Upu5CUKYtKpIw2tH53tvBDG1
E7bujhCLDbafcGM6MB7DgPOJb3eHf2gQ+eIhnUUWlF9Crv4e5dXG0C7pCuEJOHtBQkdfVNRGtsmQ
fURpsusPEQn7wqNlrgxjpjhx94jbZK3RT41yIOhJsz5LOeXF+nQXC2xtu3hEF8CMMu7cbLIh7N08
8aXJ2SnCpDivwoZH4sPMu269WOPlKuJU8WYhIz2Q1UyfzYXEJXusPLc2nHYrE/td6CDMEc+Og3P3
1KTIjWrumK5riLlcgWK2azX81hx/boFaB03t34h8rAfnt7t3v1Ka1p6eh2oqx/CekL9pP3widxZ9
tqa3kZoK/CMHnSpFIH0PAAKuiaK2kcdwBp1Ua3ch0rxv8YYxnfuDdbUu6+VVvbVEdDUbqDET5FRh
JgCjKnBQ3f+yN7Rwum3LakxTYooXsCGA3zgCocLsQuaVE0IOvgiJx8BU3iu0fMWrYUNQPR2ykNcZ
1tJCZJPx+pmvAMYWJgirotmB/Ivt+EV6+Wq6Tk1aV9EDTFBekx+JX7iUSnyFYRf3OjEBijj3bqXA
GkoWeqzHgaEaUCdvuCGUFpuSpHM7942PJw0cqBk00fP5bvqf2hIxwWqUOqc42+WJw9UP4RZOkc6Z
ZXeg+Ug7gdCBSnA2KILDjLw34NN1XW9wOONvmN5NrWJkKob8aq0NG21m6baz6FVhvZT4fUpjn0M3
rW99Z6m4IfWhPwCuX/2SSBUthIbl1E9IJqVlb/ggH9wD35kq65N5ok9MOVcdERrbgc8INaY1VsTE
nNwtqAHCbuUyyvl0mdUcPJRrG1HB8c4p/QtrUFZJnzPsiiOABMj0avC/8EJtSwrmkBpy+OatncKN
f2TsdXFCkRBd1gu05m7gNSlglZEB6ZYXGTo8dxJUnhaIluJGcGfePW6Lx2ZCJPZebNgUvjUVnFB5
Pzq0nKnYLgfB34VJjYll8pbDz62p6cOhC8UGUR+3buejd+jV7ucsC9sXmVMpMYT/aQZHS8m84Z4C
sjCI5sK/veHOOa5mN9x08kDAXKz35oY8o4/pE1qGiF8CdsBqal6KIhCoC/nin6KIQeRko9alOYFV
nEfeFqtDKsfwpMmHdSJgFMOhHfi0o+gzMxKkRcPxxWpWawmzqULc9oNzf0KO5+WkSRWirDVkC58z
kwoP+NM99mL1NkhCPNsiB4zpgFHRr0mnfIjTI6OfjXIljKFZTOcLR+oXVxhC4CCjeZUZZAGIfFLV
QL89fln3sfZEetEXFPaY2htgLRQFr56C2eMnBgczTVU8dRrm8wUoxSO4aWr1v3vulbYkZaAtcI/T
WKplXLidAZR1jhtjMTrIJI8vm3CEV6BM0YopJMdL8FrzF1qsIfq91fTGt6F5v7rjiFhPKLckoM4b
WPHQdhLt2DdpVzrTeAhMkJL0mCW8efVhlpX1s0xiEXpih5Ei4Qnc/HZwzQUieGcmn+yaXl/uskag
BT59Tuqieqt8e9wVWtukeHg/EplXUh+ZAP870BMaY1BQXan3ge7eelPkq6zr5ykwJtDaJRAptnTd
FVsI/qOKkKBoWdH9vv5UOEhUj+XQ8ugPXjiVA2l2RWrM1WzyZY/Jm2QT2q0s48toktoiH7OO9Vbu
YmoP6enxfodnvRQYC4WORC7dsDDE7RJawAMRgDeInbDsgMTbLNRuye9vG8zVxGQDiciHpCJrh5Qr
YqF7tlWMD4jEMsOkSr669hsBNX9VYhYX9QAZ4ECt4ay1xSoaxcrn1cvCVjqQeQ1uOBgSTUhdqSny
CKPOUOSiyMM0nkMaE1bt/cEFXm9Qlp6SbtHNd/ZexJzUxwGAF8CObSpKnrTy7q9X4rjGBhCRqjT0
byGXLMKRRH3yjkUuqK7yNJw6LGq27181Byq9Gk0zEBYQ1fWKCV6cTz09sr9D1H1xsnvShLs0JTvY
WvBZB0ytlTbs15A7lPZniWfKPsGY6IsN3l3OgnnezaCszMsfTvejNjm/jGSfRqZej0Vsj3ZSILAO
evr5SgvqvAcMCV14A9bl0qqeD2VG8aTaFccXRlxoxSv8UcR5mOnRTu5AFf2eBFaN8BvrJlj+vBs7
x+KiI/7fTCyc9LSC4eZsvPpbBq2yPGn1rjAsV19Gnvd1XpFJoZvdS/dgEel15waM+GUeNpxJ9zZV
eRd8B/06WfiA9e7cGb/bJXSngnGD28GrL2DKyJK7dD2z2VPss3ewXFr4ZMCIpVluLY7uNfhxBHPm
OStzDeheRbx5gDZo9bH2GgfPapfB1FjRfg4I552WEX+6haJeO+6MSZy+oE6XCFzHudFtOLMPsAnm
509K6fxIFUghd03benu0Et4/0zUiWUYRfG9WffKQkJDFSzCS88G6GtIN05ieqxJqD3F3V1aqpuCW
zqAETnniNPRQytABKjpvTwMc3jlQqOWmXPHUKgEDeNViskbiNv5GDmjxH4teQBEoVEaXwWFDbczw
4Xw+7IVyPErfUwLSkJ5oT1RmHpazxll8QLS+GDuQ426nLtNaRFxPH5NG0fP8qj1DdK8o3HX8/xHj
42Nm+DGW7HiUcPAgJH4/Gdv5JWTOJB+4b0Xtj8mIJCGCecbptDR6U5dSjkBLYJfGWdKGDGAPaK0W
UE+hfGjzt4TvUpiXCMrn8qVuAscjrFEfx4ILC5r6ZFAQiVPrhDkiudLZhxihfrVi2uXx6z3+tkop
kLELGXK58e5MHrok5vjHp7E8tTlLl0wZ0mro2qJi+QgddDTHi5FXDAr2XnJALrRmadb96EX+eTPE
nVNEzVDeH9ESapgnv5zRrjc9eRsJgQp7BRzgu6XMQfrSDSrJ+EI6ucrQUzRAD9gJMcUGBVb20YyE
3WA7lEmttx6S6O2taTJmypvye/NdoxTrsCYfB9fDSDIOpkU314FK6YQkrnud2pgZRhflaXQO4AB0
koZ74V1sxlDKzenmN2JUwACzjR9Z/JmCEgzirRWLhwmjwMcaAz8P5ud3oSwPLngqZ+3ckPebCtW/
YNd+O7AxSmnj1j7PoCCYVkMEKWVDSMcEDiUmcs3MisRllWCyn0cROPRTi1ELuS1nywv4Q792WIvK
kwRoisjWG/QhcJ7k/3e2mW6u8hgEYDSYvBLqZP+N3kZ5YbI1bKZyBPgYE1mNEeXOk81Ji2vSDhad
W0VsjprhZW1xMt1GhvRNJDghNMnoJqbQQNq1aAeKaOrQt6lQW9oInMPxjJUInXWkKTsz0YjG5YUn
fH/nSCKVIkg5CSdnbLVJWYr1pRBYzeANi9sivTtKTP7iT311gmtnzceZ72bLWmJtgszJoQSbaVIN
4Wl73B8pX/Jh+hMtTRFdb/8vT4ROkepEBP72nVFLcc6yOv8vo1wyklxx9iAGt4vdv+SAEN2XBT+N
WxFN/h/xpPPKxiPXJODFUtOLAviao0DkmKp2NJBA9W/iuYQ9Oo+aqwS1hJ1FIbFc8irc3mNr3Px0
MT13c1MTwxSlE0BfYe66aQI90G6bRle3IdAFGIRENrINK0g7J2DVtzVBEF2VSWbJ3C/2JRuI+7DT
Uag54JtGxeNF7EC4+lAHpKonS9l004upBFopRNElEcH6som6HUJ7CHA4XAVLRQhX4seIj/FAsktH
1Zercv+/Q6fZIbMPZC2mhxgZai5pLsDg00TyKqa7sz2W+yGVPiOcUD7wRp3VvEhh2d2UYDjqdzqn
4DE2CLcXvBoBe4VRKQC9C8WOXA2RiQ8gA60Go/YnXeh/19qWuCE7ICIxaRaF6zTqMlXy0RYxPye4
VujDRkrWs8xkS6pZK4gImhj1uZYiAIQfJhPMMUKoIpzb91knArubIDwRzfp0XzkfDJB0QuZYTjHj
i32HKLoyhZpeNk6ppBUp9G6ViA4FGWgdslGqRP34VWQcHqWjtAX0CNHETPCQWEtF/tRugEl4MHaa
xYvZ6e0uhGc9YuIOpTt3fGu242o+1oBMLBqpWPIQQdnxkBMNxOzVW49K2ofg2z5Bw4QnxprEhFYl
auJYvpokqpQql24QPWdCYtywkC9YLerJcZu9XJAAddkBH2QmD2B/YoQm/zqGgkcbjG/fIdT16dTn
IMFy7JORv56Tbtt0Tr5GWdBzpRk7lmJN1t1/+HGsqoeSxxXjA/ToiJX5MO4wfmGwxw6VZj39w0hg
u0h3PFrTq/oqg2nf4abekZwFQ2i3kp6QjRtSmQrMiANNSbel4n97VXKs8VeiAYoUlhswqPIzdpmv
TpZe4hvsOjMJBszz2QbVXxQP4+0KfhwuYMoSPsimvuvchUZCsInSNuIby2LvjXlfQUjAT/DReEL4
mLgRqqL50Zs62negA+URRrmx5+0pzJIZ99tUI54K9HDzatSYNDqnT+7BlqCbHUWQPeodESNd8B64
aRe5fcuYTD0RUDu1UshCjyYJCRErzeD3xISZ5lAUqgdew7GLsmz/7NpX1VZSdk022VrMbBFlEa2J
xBn9e0853q3IDj/e1d18rtruuU3bxKSvuk3fq4T/ay+p8kWS4EP8GN9TxSMfSFp4hbrKU0J2gHC+
INiexc3GsXc05KVir8Ku3CRF913z/WAyWO8THulZtQK+tsEglfZF3oB6XEwq6uFEniUBXyML2hPH
TZomzdDFcWiF8ArZ7EQSYmZ+y4AqangWwrJoqs+Nn3Vb0Qu75XdW8+ZnqWuAH9fr7A8A/HvWVwip
s4gfTHj9AhRhvRwUwHOD7xJyAXDW8LXC7FAw7i1gQpOAthoL+WEnzGLukhZJaWNcsql2R1RzzrvH
EWqiE/xLZPmPQ9+eji2128j9FnZCMWU+c9xTjSQ04qpbVrEiKuzEYv0D7E9sKH+WKKh8bxR9u4w1
2sxcgun/f0gzuawyMmsAfB1YhmSmUQKVcgwEAm+EUgF7F4k/upVatFCyp2Bb2XpmCIZOfeVF1jLn
UZ30JaM7RMX6Uxcs0Ms83V2pfz+d7UNwhJcsV2+z7VP5ox00n8l8/3QLHTPcVEllIXLPMAlu2epr
iWZyL7rI1UltIMNNAa6adnGQi2u5vI2skl/TIOgwJpJii/NLEJCGuDEVujSPc7vfzLIK4+CGZSH8
dvDcmXPzSm/M8Pk2gkrXZPrfX8QSu6VSi8w2tZGwunyXDZDYJZoMNis95li1EOLK1C1sacQDae2Q
/dBD97c6a+2cCpiPjCr5dl/cvQlFOwLKuVGAKHLDVhxk1eAn2oHH2XGRUq/ZEzEQrpFOTDWnzzmM
z/v8WDiIovZSRr4kcwO9gKQYUTTTKPc5DWuK1mkA+DyjB4LH9OOaSh6njv4Qb9c4RwcWQ6RkTnrV
rbfujEWS9xDZZ1lRgxzJj5UFKR0JonmnWT3jr60Qf+wpHEeJShXNPDg7AQA4G4wtQw/qFAFrS8pw
EBH6NHU3ZXyz0gsP9+e0+Xr6Gr+v5bkatjjGu+PrT+2oz5M2bjP9l2P1PKTrM168Bq+UH1ZV09b3
C3wwYh6Nkf+zpxqufxn4GPNk512ppOC8vMLS4ULng1NLtmRmFsq3i3C4am4ejd/3A2OWgxu/A3/L
NOlC/FumSoqLhnX7/LRKSkqmAvsLUHJ7JgoN3jFzqBA9LxePw+x/0Tsttj62DMLCjqXajWn1jrQO
qf4Nqret59Y/im5h3MYWjzEI7H8Mcxg/wgB7TaGQ0kSX+BTo7epNzj3t9+GdDSjWX03mlzCMcbT0
9K/jv05bOsOJAUwUHg63jTMGzLzZj6fvetXzwl8v49+NAjB/X7DgcYeq3wv/6JSFKMx/AJGLTkzN
ZPXSkNnbAM/ISO60EfMeeXljz8jtRmFdceqLsFd4lqLsSdJWP1SsHXeyRH5XTppZ0YALffCm/k+g
GGqBRDicrBV4uT0z1hbSVwXAM0qj02peQpELBbTzOkkZHFsdeuOOfbF22BQTjyu0WkM3cmvONv1T
UL+5GDnSrahK8kIJxIarCKkdGRjLzUZhCfK+EXo1ry7EEYci5lnazjMRXuUqgm6T22ryMdJ38miw
hsZeh2ZS0YB09yiguoMblnTQ3opxTitOAi+eWE1jVzndgKKfARzgjr18aVYQwqvabsJY25JQ03RX
r3oawveXsFgji+DY64Eo84VXzkXOKtu/tZuSkDGH0CXWHW3ZpJfnI0dop87IXCHl0aKhq30q803y
yJcg+KYzktaBLh+sHzBWYhdaeOcy3nARkdcRlu62KAirvxAMlkw3nLwLYVEZHYYtDdiYLQOc5lAS
d3h3pHC4ds+7hrwJ7HDIhEHES8fL6hYCd0OMQ3Gwx72BoksRQUVIEXKdpPlW7JmIvikX1QfXytJR
mButCE/S6t2X7Bso7+TLJgUASoM1sEqhvs/ACFq1QdbaPCBTZrstlLzxbKYJKzIVLSfuTHxCbwnU
6Ps+BI24HViq7iWj8Q8eqKxDU+VuJ6XzRsv1cyJMq0gezghw3qFcnfKsGniDRXwBrdNxtR7jL3Ty
IWHFxZqdSEvL5I2aFH2XhtkOu+UcYHSVIW5iijT4I5FyewiGtBHMfn/HHaFnV+Sm/HpkeQArqvD9
kGYSweoOiZ9/R8iWhF2GcKsL5fpHZ0NDgMbOjYumBPUkTcraT2wk/ASw4tHOD2Jx3zgCUIAFMDn/
AkmMe4aNXd/6WfyNyWOaHg0QIkc4ewh8UiFMRrOwLoTlaLpLG3k1r+VG11xp3xBvXSehPe3rw6LM
75biT3iohdhD13dWry8wB9hwQBCho3m4EDOGcEyc9AlI9pE2YsiRU2m8MCDzrmnmrKUT9EnJtyV6
QTcL9fUtNTod01ZQALtR759ly2hUAU1vSJny4A4f7bR88cmSj0V45MY5srUhd3J9S60enorFRBes
+M1vlooceJnZp2WOv1NpkjhJCbuA1+z0UvbIDBzC8DBKeLfgsXnmk69ObvJzfmZxMMwqB/yNkoQL
GsAGUj8L25kx4IvPMysbjjhZ7VjTsr1Wv6wWtR5pVh0aDwVQbWJFldFuZB1AwH7wyMEnHRuqYtQz
e+NpFKsK4FxfPDffi7k0nguZf9sSUVzkLEhassOBvzDL8iPutvCzEyn57ruUh17MTHujRcqaISbd
HkLKGfpvIosZQeukw/hNIn4oGdHvHse/7EKwAkNvMof+We5ehHTCi0zFqE/z+ihKidYShW0UfY//
QsHJUWmphoJXY60kelVJunZ9x4tRdwyDFOU8cMQkZDX+6ITXDFaeNhOoPOH65GvZhtmvdb3nO+xa
obUeHlEeuUPhUCUEWK/f/ZQBRcoUChc0U0qBvx/goFIFgbpkx1I+ZgTAx9C40qUC+mPAggbqnFww
h3FrgxIQ/kkxTsKRya4dTPnYZ4kX5cF3mxeC7bRKe76WYgLN3RgzSTcXQo7L1otEUa6e3tcZx0gs
wojdeXaUH6Yzgw9jpG0usCPC2twc0KpJDMXN3ZPpfYbPP2qNTYYCgPkYlxCr0wDXtjb3tAwRqTE9
7kB02hI1uTYYUsYMblzQiMBDfv+I0m9j2DJyw/VZ8KLubR0KKz1DiM/DXtmYt6i3v/tNkYsADt/d
L8PQLA6n2kHaPggWW5+eot4oO9rNYU6QmMkEwhyp6pgcqAJmhDaPBUF0w8JQgLkVLWq1t8ueCrs+
14eVWKwu5o6D8/tnxIrnKEVDP3G4J3OUwf4XmN1zXgtaNljawwhgTyjgH1EMPtoIZdFupyg7zNDC
bt2XcdxSHm1Ml+Rw9ehjQD7zctJClRJbB171LLOwDdqqsfE0jOUX95usg+0FrG0t/FsnRoudwdeQ
mF/PvjSqfhwMTadcPP7oCMjN9vBJNJrDYWI9UpUj4KxBUzKS/07UUoJp5TcjNEdm/jhrOC0+3H9S
ghu44UxiDN5H/ROpPgchXAmBErEwgV7gNGXtdsrcQCPar/pOwyicEaaG66YdZbDkquJUjFUtdAp0
daYXKUhUOClWX7jEd/IQ0qKDQucQzPI4/9SJFr3dyOXEWjc5ECi1SpP/tzW1spEzrGHYtnjJQ8ut
v4vrL8vn94UHx/JyJ4nMvrWHGjbThx/z1t/cmHHhI7nNGZeLLQEnZn86MbFLr8suYPN7bSLFnW3f
F3i6qGU4Hjzdq4N/bc+sI9cx2Rlb2Y/PiaXxt1fQz85hJqkiFGVpTFUfIW1wk8jH4ipQKs84lRpD
6MzcZNkuwcDJd9PRTIB4bFlkOsFRgWDBe1S642gCWmNvHxj/VYVtBQIo/EeZ3Qe4r0bI31h/hMMJ
vm7s/CFeK1W1YxUenkjl8IUdbJu19DnlWoQLodSdzIdpAvqRzGsvDUv4sB3QuEvhpDBbUfIMIeRG
vtwOHmH58CVl5y3qj8+sbvoFYAUv/8aieP4vsLmTCLeBP2pKydasPGnnSzmMADWVH9Rh7aGa1ZUI
QNIDysx8AJ/L2AQojJcV40wgpMch5kiSPs5UfEGCKJVQywSHdoQw5rA4SCmn/Uyuyv11ivDYBsx6
SzK2Eu3Qf3k/1KJh2Zne0RRAc0qzjnf+O2Tya5nl5QdKbl3O8WauZRkYoL46LOsjsVu2R8yz4Tmr
7WaMDkx60z9LybZU1bvnLjnlpa3gUyLGOO+ARlbMtdzlA9kP0XyiJP37Hq7NCZwq00c/ZtGyLloQ
BGTEn5w5WwpeDRxrJrZ4xEgr/JdeInBKSWpEjDA8c1dkSNisycsUHzEm6lW9e0mFZXS/HfqEiAJ1
sEhkIngQJYg8gpl7TOIdYNSX4nOthnhlCqmgliR7RNZLxHYuQRp+agqbd0Jq37SqM0XnUVz02zBy
t7kM4T+1aQmvjUv+JiigJa8wTDCJ4hu/+JbIzXhNRhf5ZZX7SkcC4b2K+DPicvneGDrW/mmaiKWQ
dtVc/MA4+3qAsAMwiqvQG6OkSIYQuciznT7oI2Xmr7KloUQdYguEsS1mKOaUJevChMx9ZTlVJ8vM
5qGA/OgiJX1JulfJwz1hX+Y2NxvVGSo91xsN/Dg3D80u0pGcMnQhE1W0R1uRPpoUHgn06u6md53W
HSJ8cPkWtPdnWIfJGckr0X4wv5mV4NVBuKA5Wsqv9QcXOamaDjf1XlZwv5nr8zn+aHnkzw7n/j3y
HntCG2o+4wa4C0ucxoAUHg9ouwpVQB3tvkSK/e/aX7M0GgCNVPeVhENiOybf/hMrmBoysYFQ65nQ
7ag6QB+gLdTLeD4fDaVzzoJQtdnPnvcGSf9dMBVrM95gAC2bgCw7W4Grqo1BmmZM+X5jcEAJs2NU
XxxnShZsGT8EtEow9DCXiW1lDnM1MGP+DMvpkAvgHAV7A0nR7eGq7MlOI/O5j22/LJUWakA+1EZu
FVvjcnjvyfZVIt9MyZLf1gn28hP+j4kEqAJItMro21962DfoV3sbT8+eVZizN4b/aK4LMFpqDgVx
6fuSc1CF/V8CdCXs+torn/BQ0vmag4ZiDQMVw7waz/1CxtIq6LJ6DeqVG/tEpR68Woi9kGsYq3B2
h4Mk1mkWnMAO8QeO5s1oEL6idf1TIuY5cG1TU3kU00VHJfCnm9D3QHWIo3jf5KwWo3492H4ODISW
vKsIyV5FzOoquJkZTYsHaXoGDGpI04uQTubvSgkv60Lckd36sMn7OnsQs+EP3bNEdblod10Fhe20
bvPdAxzw7o4ZHi6zoi4H2dbpZsiguzXJQI7srfUSXQ4nUp7CXtilqEoNFvvGsIB6PIp39/XCnkqp
uvm62VFc+2GNLIYWe8iFMqLoYR4YUtXThrVs/b7eytZxrm5uTVyKQHGaJNBr9Tos1hMGcZTDC/S4
KXVxdDiaAOPDe7I5aMDw1wpyyVd2QCsHi4rp7doJIODAwTMVIp5LDEfGFSX+RhwBrjoZXuoomm/b
57koHOqBI3VAJapI0eerifillrLGllRbH88kd8XfeAn+AA72zzmbPQs4gS9kZrGhON9rCsRtrHJH
8Hwg5yg+It4zSAbSXmVqdGMU54SFKPV9fmeGGDvtQ7CYH/BUo1yF20llkvSfZZgUhh8VINUo1m3J
Rk6/EKJAB+cTzPFCuvbZicEqMKe1AIEKHXkHO8C9JtUUgqWfrTvrjISaJvyIPRjma9s3wBWYA5Zu
iONOnJpPC66ti58/DrgCWYuvBwy7zblFOsslB2R5t2xZTx37rgrUvMpEMJBMwTHRgDDVS/L/+XMi
xly6qcsIsb+JvTnp3mzy+v2op2d6Inltwy4GLLQ5atLNeljutnJb9EbzBkRWhB2A7RKyVDeSN+OG
PVQkBN1GpBLhZJ9ufmqiL4ALm51OlgHpYVRR/RiGE6kza9R+HFl0MuIwfbs7T7fRFADvEW2c1oHn
z/SIdf5YUxU3QluFDeslJBcH5HUYevIXSvsfsw2ozqSqYV+AxqexmEiM24L0B30eQupGXXE5hCK3
8DJMmQvQY4jTwKfI4V3t0lSwT4/7ySX5f0VEC6RVL5HEgOI12AoM9WHNaqJu5Y+YHgUNE1uH/MqB
DjFHNvFQ3qQBaNPdGTtrL51M7Tgw+9ubKRsHAm5D5ndxqcdiwdlxY3Aa+KE3Z5AS0rVD3kK9NgkP
97SCRbv3EDb86my14c/uIBkDkEHBf1z4DD/GS569fMMIgu/YrvomZ63vlxfWZToGUx0mcM+4Qa4/
HmFbrc73tN+6b8P/yIJv15Bz3wYodPQX0lf7Tfu/Yh3Er5lVIwyCY5PHCyvXHze8cLFRpfREcwef
MzXA2XHqgaLCXSI+WKUyhTONIsYqmofzHp9i3KUWuqlrZ9m86Iav3uWZaKMzuqy5pgRycSPjEbiI
4XjfrmXyRxxe7ZDZ1UljO3WapQ6u9Wk+PzjBxPfVzmTt7DM1GfEZB20tq2jElYZp3a6VaPSoNwE/
za5TVmwmXWaVEuzQljOjLOvGMo+a+spnKddYO9lfimQr4OH5b765XbH2nYeuv3AlKw9nX2ponmNd
rkqplcmgV58bHutwc35diVjDTpNl4wagguuaocNZoDOmYrAFX5g4F9g4WP+SDolpq2dFr2YDn5kY
XzykD/+H6XUtsGY0g43B3obFcfpCDZfMaoTskkJsVkD1DF1HCr0IZTh4aed3CWXMYqG21TDYb4Il
ssjAv0ykS2ayVnTM81mz+dr29LMxMTPjwjfcmYCkr3DAd4Y6Oe5cpjmBUiJglUGYGZ3G1Q0i6vwM
5Bvqb30GEPetIp64rQ3YZrPYfy42N5O3z0tzy3vdHgpqVVzEkWm4cuLx6M4DZtOSkjoxyvDTVpG0
qn1CJHr16ACabouZIY8nTXcVR61ogTTBBB/n+mUz2/M2n8sJeJR/0dQFoNqAzUSoXA29cudVfj0i
3zTwcKDtYUXCS7mOkghphIsdcRwX20vVAl5UF66fhY+wwNo1hA0RQ5LaAAjTJTyChOQUoM3+/+YM
Vl+IkSY9EOB0qXOL4mT83Z0tNGzAQ8jPUqxkJh/p8ZTKhKEIYmDsFxRrLwYBwKeaMdZKrjDJCV6E
AF/svWunLoRgsuL3M5g1SaMVUSTetR9eGTJJMBUZgNt6XYIDkbP1AQEB3JhnNtb3mjdE02zCwK8/
g2yOLDK9fLKJc1gmKHrBCD9BQqunf7jzqKMaKiOrie8dSQFw9JoN6NnL+6BHgt6P1VaRucrlBfDr
0XXY8GFLONH6VLEXGL32nAxTbMkxoxeeLIG9F/ayT20/E/cyMQ2N4c7JSAK5xbf5MQicijFxAPFZ
DijCqgxpICPfae/7LGXR0FJbyILlls/0hQFwdjFz9PD5BHTKGEAc0w/he+O0A2U7VyR7Bh2VW8AK
qNhy29JNquvabgC+ANhLIRh8nVYUkyhgsT+hx3xgJYnUn2V2aUQH4onm5eBtCaRF1mY66IuTmhL/
t+4JecD+xH2lqkKwfApSVIglZH/63G2YmcsMFT5czU4n5aSHZjIW2vvk+LI9bfYyO2Jmi73B7DRH
DENq0UryhEKPnd8B7GarXa9TSLx98EEaHxRfuyUuk16Ap2m5i8GJfTgI39wimpPn1+lwyw/P1ETy
bMHqW3gdFSXbuP1LLi6ACfV+Keayoxff8ojs+NjB4u3u54nOVnaSuw+6BbhC8uRbW+4xHnUsf6lQ
ITX01DA+cjtZUkWdg1wz4EYXVHXq30t9EX3hyy8pJPiR4c/JzgYmKP41WdmcFNhsltaYaEr2rQtL
XNVK1ILcoFPpvV/rdVXJ8a5sEQqxN6xpGsBOIO8FN9mJux/DV+o3KRcCP+Fm+7qNGXiO8qfdM+lz
zhirOenFS/7iBltH/JhRe5qFQ7eLAk1YhuWQk2MJHeuOFI5t5lNrKpiUBurApbx4inNBmTTOWZF0
5cFJVJ/Qh16kqhY8A5JAyTlhPYwoNY1hmsYQt8pHuTO2hA+FnBclRTjKXwxiAVQNHDUoHiSz/NgU
UNYhMgQS5LCHxbDriwz53kYeS4YHGd7jW20aw6Iar/5ketLEUQHnqTgs/ToYYpfE+iKaXlwrk6DA
ewnStBzJ+jHf07XAH+0G8+LVPoG3DNJJAGTmCJhTQN69/p7oAk6uMRoqfmmeDCjL9fxIX2I0h6dA
4Y86WrSSf/6cC1d6gxbM1KoE4SySR4pt6g9Zhvhw3K2browKhn2AIYkGWnCbKrSBccGMp3Z0q1Qv
WZUTajc4fCGqW+HdqCx7Mn7EWYaTc+xiSbTsCii6LdC/22U1S6QbrhxigXNz5tTQAeuWeZAtEjfx
fxbiJMu1noasKgmDKblKMZH14mRV9cJiMvD7zq5tdyf8sPCl4InfcwNDGlu9mymodnbEtr5JocrU
IGsMQ4z/J2t5TBb8Fe8sfY21ON5v6yq1PXyLFcp2YpWuerBwbhwNacMKEukZFHmZLAxgP1Suh8Q2
oyqVuI2RH1TnSHvpXJQWojFWMH/x6soObl09w4Sh1IiF3wBBItJV+Vl3Jx22rOHPgPsEp5T4x54L
hjmV2BHoc89/J9L8TjeGTnebTYjgEEJM4Ac2iHLL4oK/ZIGToZtRBNgqAHmaNxX5kzojCD+9snzH
nyBm1N3aSIBDnql4lG1MTciC/3dMs6mjqaz4prnGBWUKTjfAmXModNZB3wvNf4kIyMm6apYWoXql
keWuwKeIu1j8Hs7K9547vX54EWyafCuvryb1GQAxyHZ5oZIXAwsJ9VoE1gN+VgBcRY89YMo5ckd4
fEBkL8gW3NN3BmXKLl7WZpudBE8ZG5P2U3m9uFLryMJ8gNJbI+igIIIdaQ5cqIeOl/0fuv0XBUzO
UCc3/dqiejoBZoTd4heqXXktsu00/ks07V5brl1OPzEvvU4vyJdFcHG3xbcEhauQXB3VaIKKr4NR
cMimc/JFaXVJPE+T5fiBHfP62VpJ5iIPjkW5ZPSzmDnW7hQ3eoe/gbNSLhSVH3zf3NuoNalFON13
lDkVVAnM+y2omMPdlY4lLpt0xBM3p34MpGOiGcsd4LhOSQSXqYvemuUEQfNt+PBPeRQYcX/TCP3A
csPmCGyF8qq2/ZArdv3Kbj3AmlKFKlamHzHEr3CkIj14nSLKmHiCrdmHKsVS5Mxc29ni5MWfFB9d
WbB22loLBJBysCoNGSyPV4yoFoX7Mm+etNOrvGLFFxQsSag4AJeIjAlMJQ6Crk0+eyOVsPjG67Ub
7b9B77eL4dsLNu1V0xeJQW7Fmdkbb+VzLff3x6Z2CVkecqUSGCPmFMTbCl+pWJFuWmfPu4EqE+B/
wTWFKrjlKdj9dfgnzMlk7wCub8ykkFWXjluyQ0C2EV7jqp9R8B75LzkS7ZGt+94yrAMRjFMhYPTf
1ivrUijGA7gmctCtR0wciv0dxayPl/fXLnxKhbD9X9LBODaEeSlN1vQTaND2CwQvlWZc7z8lgilS
414xnC+zE7wKXVKOD7qOqmPC/9rUZQx7Rf2QpTil4e7CCVbfdBixT74dmo9LI+/LVZYtRrszi9hA
6HCDQqf8/fDp6mlnPKWEF5XbrhBtMzwBydxew0/HCfZF95ZVWJIfxGPJx12/l/T9YD3WNGYlR+S7
oV1OWVxSu5rUBxjsWjd9Rof9Y6GVjBuccfBjHT4hDU44wdKDWOzd8X3BwzTGgTPn8Eh91vcDAe9o
W0XoTTd8VXNO2FACdLYteMw9nEYeRqUX/7I/iEitFy4gfE/YUiuLranzKcE6UqKCmdtnqLGCUvHo
ERAKgbUp5uXBDzQyXqrgb581mgh8PzojEbw5Sl0DfO6J9wn5QWStc2poLvCwU5ZUAKJij6A7UFCl
k/PusYuHjLt1uqhmZ+E3RY5+Jw3L7BN8Ig5Ra+Rgs4lA6jSOP2kN8+MR9xxpclg8Oj0Fflam/A8V
cUJYOXGxUP69M0zI7XQenKWN8yhN8L0g9fiqtLQe6XDtRR6Mcwop0YP1VcA3b1hnj6LdKFWsgcDb
ETvfXtT6bultPfMdiE/lTPsRT5xiviA+vbQb6cc9FVYzXHJ9zsE7FxwNCTftbIyuBiupaaOLMoyZ
bTxr3XR8VrUYEGwmdATnDG7GMosGqXlsDhGd6CND6hpXVIiyGw6faq6La7Aj4Pgve2v0K9XBCJKC
HDrexIssucQEjkasUSzVvuYvdvNczy/idj63Xjzzu3khYoQpJlI+XUAOmmiPFo+BNuEX9cl8LWJM
gwGo/CCZ/l1/q7kucaXhUEdHb/NYt2d9JasbjtPnBin2EHPa5QXyWdsIup1fGJAYxVpHFQjcU118
WoVvUbJACp/yrbjoYYgWxMB6Hwd4kHip78nZE0zwASNnDfUjDpqILTiyWYK+3VKKssd5r8oPJBVY
k/hovDEffAAUQNmlKGHznHQT1gBbH6knSpO0BQGkbdn/IaCgaX0drGnRwSfLME4PchCUmiAuLiot
lBim1ZZgEMGAhMSy700UEnn1byjSfjJMtiwV40y7DP150aY0Jz9oG98BFGB5a0U6Buyd83iXx/2h
gQ+EWxfHRSLB4XXh9q0JVXjwVgKIqXuljc59OByXdJsTuKRa/NEnx9nd+fKHQHmepAjnj0vrvV+f
jQhadDQ2OKqJnnK9tvLOLvhdi+ru77R0d9bw3RZifpHCuDdjqwmu+qsHFrGvurKhm5BiLPzix/vl
+wgkDKAt/yx+v4dqPmf6vyxyg+IdqqJNEzrjAFjhvudDm2ErucRqOhN3dClRv1n2Pa0C6QfnC2aG
P053WsM4xMuHOyUxrEN0DNV6WyLweyihKkqlXb1snlk5c9PuXOLdpmTkMCvL8284fCN+hiOrA0mg
aXtyRT3lFHHlM76lS3+Bib5NLoHcC7km07efm1GMWwQBrW/oev+RbSUCZYE5lLJWcCGm2/NrfAjB
e76KiX94RJ41x+xhKKjejYx/D4QQAjUf923e6n5fPxr4Nq1TJ+2S9SkIvdn3mn7O01+nxP7UV4HE
isJXW5EO2NxX7CkrmLP7Q1XUguS1KXL7bd9bJiXtjclIq6J6fIDOy1MaUdWJUXwFWyz+MqRkbpN/
Godun4VDMDn3Np/OMamGpqEfnt+N118+Lx0jsVWDkiqA//ECq5ncf4Pc6W37DjDkWVh8Lkmg9KXf
G5myf40HqubwNUV5n4u9ot/JueD/C+IIROhr167bMYz7SUS6COwpuG7PHa+iKDoxbZqQzdNFMbMv
Qn3YGy1BQqqAWm0/HB1xsU9+sCrelQZbKLdVxCRpC5xTjthwrDKoPMTRaDSfyAzH9lxVdM8lyJjF
HFtjnr7HlsDBxqhLb13iCfNCTRzJazX+U0Pv0TcXWvZ6iwYjRE0zdbBGJ12t3s0WzQfFJOxHEqYl
VBTk7SnLGz0WZTf+A0OSj9oEcmbEFRb2pwagwNNu+gp5yiquoGmIhyn3DR/QsCa8tlDuNwqQdUBm
sRcpuFOTqQg4ULdBIfa1dlD0E3W70xSJu+qOsPrLKerG6q9ILFakXL3N4O5iUC4c9TOgKsQyerYu
B06XkcMx8/aPBenf4pa/V3IC51n0EOuv9EKv0+KynK6eprAcPPVJ82V+cWdeTcOv9x1ZOKrJSw4A
xTyzoTU9qpdmJFDfsrt+gH2qPt9w9CKj2thtNS/FNoNhTc69yf28YdyYjXgUCw29mYJs530a462n
YFAM8KIScd2EqXJrXw8OEMoe6AlF5wCDWQoylTdTGLDtA8s1Dx8Zn6hBbqpRMLiNFYFSO97ur8n2
99UFco7+3vfLuQK5Rvyqz43rPHQeDtBQc0hfhWIqrCSzuUnNWmwweh+cin9M4yL7763sMhHKWJ0q
ZvYes9C4BdakiFq0AXcV8dJ5EfbHOxMbN/6+WLb+gA+Cu2mnQB92g6CK5VgcVW2+i5nR59RE/Tfp
O0hRhOzFdTSYqCgGUAIzBqxZlEo43LI6rrsJT0H5h5lRrF23fsPKHRnJTjOxuYAWvyERhBK74szf
0QU0tSBgEEjff2tWVHZetG1b2bXm+8jGR7Z75rIQKmwnG/Y+jiA5BcTKG3DAbXh5RUAhWzfCJz+0
JtwPF12StxX/xBZrXYSQNLQ9Or6KQ/aKPpJY3OuaisHdo8mOOZv36hxQedDgqOq48yLQwLsFattg
28G/1vLdA3eI87HQi9Hv2ToshGloBZGt9AHzNJVRX+DR2f4cYyi5HNN0qfVALue9zVFWgBsolRVq
lfhT7qrG2h/PGkNAIjmOXY/P7FKIk9VrfzfuMddjkszsUqQ2A2QKgCvvOHgxodo8aDoA/rWl17cr
ickI+vNMlDQx1XnH+/kQeAamQFSkpaDp8j0cdfveLcUNDrm0a7pcIvX/923yyK/UEXcYBbosD1tk
21fxQCjFdROP8kroVsBLwSyKLs1TQ6VaNQiDtnrOUNF+Z7RtA4t9y49xDFtTeFOsnz3BSYfgIV9V
j3AHHFsHfc6VTWB8YetkGW3bTG/ohd5U3jjRS/Zpjy5ujZMTDKLOPTxzzVm73ARrKSjQumaY40bd
d3UtlIlyFgfMq7KTE/KoAOPIha12HjGC65L8pPrxV7XbLYpCsTZBpu1L8c1195qzUjZdvkY7FnqU
fhon1sy3PwIT+LgTgRMIZ0B3tVj2X8ozUCJ3qR80ggdKsDMW/ZllyVRLuOnb2su25yLHnY3xONIB
I6HpLcR578d/a1AcbIrft9JC1waj7bTAD9wQxLIz2vPn/o9gyDbZKhKAe/WdVDcvIyibT8RSgh2a
XYIpB5+VLUGLjGecld13GRqhLUUnhznqWiwqoQP0CDD8z1A8uoL8wBTv6xzJanO5Xyykstx8WP+E
aDdXYD7e2wM8iIBFvt7D1zlh/MR/O373Y6rM6GubEshna85XjA735GEOYFXrFEELVeirMltXRVzm
OhMb8Me7CcKBYNtVH0j3rMO9tKKUJ852AiUKuBODGsYD5CXcmDhT6JVRbHjDkAYw5QEBvuNhHlat
wsyrT300OjF4qlbxtgAHfoFTSrG4sg2EFeVUGwKweYW8zKOd3hXnCrc+Ckw1a/jY3fOMCCYp92JB
plabPtRVk/pYS1tb1DQicNAUPuMksS4bFQGQZBc4nxp+wB747D5e7gSS+zjb7YXAjliAefcxTG0y
eHzyjULT0tBvOur+KvOjgHLGhiZHVs00luz4cVbvW5dx9aWqoJAyUw/lzQSkAhtQcqzMrXiAQNEi
zgqTF2rL8Ah62nxpLnBxZV6EJdaV1LvpNyqa/o5+zRDLQMXjJp2iIxlYG3qYbd75mqRdx73Fp+9x
V71fZ7kFfisALFs1LQYVvjq4Z2IoWCgRjbBZT/p7LfZfT8SV893dhRnwjrZpAqExrKETLxjhWYYh
eTRNN6aC94VnZFsiyqHnAoos1M6yF1hGAfXIkTK1wR11AnIUYsI8q0dq7xy6CwHPaC/O3MAenKbj
dUH0BrTYOeTd/NLJ1zLDDLTzTvNAO7BU7dLzG+i1PnKDLl84ByyPW6nUyBz+ZNFAVdqF5KrKJ6Tg
1PCiWK2ROtnG7Nw1Y7W0DLuWnrENFERw5TfESKfs3WOF5hTxmEYGxXLiZEvbbSquZ3k/NwNyqic+
YRmJnvnzfZdSmHmLs8gh+Oc80ZfF3D6ER5hpCfy4qx7XnUdgEFLJHfwNgbEsZYUfxlcMnQYg9C3d
XivoWANuy2JC9ynvXKPZkgyIDeI3rdhYXmdw3HDIJWclRiSFdBq+DU5q8B7/0JRom+VMU+scCGmo
Q3pv2FNrB+mU/rD+mq6UkKgWQv3tICQVdPLrvsKwqJenrCFwTaupvGfZYrdxT6Jjx4NQXGwtSqXJ
9AWSRePNaq7LkbbbJIjTgwPguMi3XDAB22/53wwDehpseoTTU84VUFVh7+ftm4+5QZqy1KgOiPcQ
0oXyxPCkBwVj6DVXEOn49ToBVXkamD0TGPjYz1OnNgUFVtTp1dTMBIpwSH6zGnNNN2bqLvU6pmN6
8MtRw1nbCa5ft7c3+qsRSRRiL1Vo7gWhNOAzgn0JfaUDg3GsZW+LbsUpcEdERSIi8zBe3XLaVV+2
cifIz+wcPJcwbmgKkO7K7+oN2VLxhETdDJIqtPnPmN/QXs/rpphv3z7r1UNdUsQzYnn5rHZdyPi+
u+q0Z1zxt3M058NCZRF1bnHKq6V93JKT+pe/UTYRWfXSHkJzg3hZiKFzSHgfgI7WcK/cB4Ba1/x4
H+nPVDtaa6jqqkO5IVVg1P5cpuykGW8bQWzeJdBil6xv44uwH4FMya+ptQP2hkhCvgu/TwNmUE/g
jnhJJt9xHe1mBek289VlTpgd7b1qGsgBj2zGoyP6h6+L99n2Bnwyd2kuENTq6SW05YV4/E/uwTlM
GmZqC2KZ3jcvCZnVFerN1yPkrg1DgDZvWhK5gFSWRx6nC9OIb/WLkQjZJDi03x697GxhiSOhoc9P
VyeaV4bH6OM3oN91E4hcSHDVhEDNAAmTaonuK2Ksy+jr8hXtgGTERF99+xuHnGF9akqrcujfDEvZ
ZCiZAJpqqo5pDxWyzPPvqf6jwm4Pklthfbhx6PWLXbTfI7RHEeOHxHujTQB2l3QFv0USG4fDANgy
EEU04R0JCC81+4vxRV7GtOxXbgWm7pZznsNAVKrrmu59LmVzeBERL8jWzxMEpD6OAhfTLrnJJqKu
RFdBR9wntes7Oo0dg9ls38ygTigrC9W7mL5977mW/BW+IbbBtJGiQ+Vd6A01fqTLQ1xOyNWNNCZE
hx+G1vbtV1r7PNNdWeAqfNzhuXUNAgrr19pZo6rEkAXPqZ0MRSrviKjojY6bNywO0HCZ1x9yKDea
qz0lyktPl27q3UfTuM4cjd2bJX5Hacd9nkUV+2oDd5nx34HdVXxBTNHfx2T/BvGRj0xbnsc9Woim
tAdrXRiVABfxdnrLCNBsZ+WvuPyGKAVYTq1+uhIfsm8Ffl1DDJCRvOreYfBUjRAD7+zMgL2ppaaM
raTwe1P/ESnNFE7NZDimT+DfsmK5++WIxp6j3t2azBrryxxTHGTLhJW5vDYL+8UxaKP5QAL/Oy1O
srk4NUubXm1pp4JYxh7feSGWaqbGRuNVNhL2Ckc0QWsaSKWmYcMlb+YohoWpTS6jJsgmD2Qcm42o
r9O8ohXJTe2aNb5qOnOXqyE6Sumw4nHKdie620pvcWOXjH1CLwXNdWZ5gEmD0454MTALbDGkzbVZ
/lFsvf7xJ+0cJrNjoigwMqkFR1z5OSa93Wp0bX4zlGc6pTUeQJjLygQNoA2ahqb1hSxbwInjFAz+
9mOAqBsZtpW00IN5LrrnkYTEYWk1rMSXmWPb9jeLlG1TFbClOpggQqnFnaNTLPkMNSP268i71q3r
7trm7RD9WsDX+Fo+mn4q2k/9sm1cSAIuxTqXIoIiShcPlj2DSGiIZ9YIE/48Xg8n7W4r3NXvkxnY
ktVIl01yHPftYerfWHFb4nMYJnA0GqVQOpUY2oir1BHal14aVPwPTBMpQsvNFuvbLjKor3FX5Vwk
9IA8yT0JTpa45B5iH4mjocMrn6pQqmkhaDxCvdtFRZFIk3iEBp4T5WeFCjE5bvnWwpgT9pMY+c6E
sSccXykEEemcDpHDRZChS6An2CPpZoiVjDKRPI3GL7eOzoJvDJLF4I+iDZAwzgt+JMddnECfKdNx
v3tDg4wRD5NbPXaBQ6Pg6GFSB2t4f9Un394Xb3xPbXg+wtb7BUsrYgMdn+v+bqf9n/5isd1KKj8l
PA6jH2aMx+aOAvhpHVhRiYvxYH0UBkMnapQvEtluWZA556OU1NEPmQjth9UMnPHOmNB2Tn0fbAXU
32RjU6qleJXEo4Yi/tm7ZJUhko+XnqdySOnKjA22gzYkUBXjC+DOS0N6Pw0bocDmCRgPidqrGOjY
AgpJD/tyKg3gkpFAgcDSESw98t2kWKHOc7E23Bj1qZcdVSpQ/qZSWsDGZl2c+T6Akr9oiQMQUANZ
00be1SV4VEbXO0L6SWzpCxA2YXe/62O72N/7/uAX5Sro8CVZfEHrOlBIbiwv2I+WMeawrPKwoE9T
8cke9d7ThDFcJS8gNJ2J0TqkaJiL7UWtPfVLtFRUbWYtUxQtPmwJsNTH9SeKLKFGspXMRmjS82oN
IlPzC5GYd3Sw3LD5cx9p9LQQocWeSavFMqUnzNMdaBDG+fNiYy3tMlRS9i+rabvTB9L3cKyd2GLs
f88MXNE0YyUsQ+/2z8Yfj1nQ8tjLmG0XtlK1LhaFW2X8EQvfghqLVJA+agC78i+g/VGc/MseOFE7
RwwvcjIYAEoc3lkvpOHRJlSxJyx33oLm1mgzb6Pmd2XUsAZA4DeEfh4WNMeycHB/d+onGdrj6i+C
6CBHrxNbup/fUwyVsjFb0SLStfpVHkYMarOxpvlod68HD45c9u96Njl9rJJJjrcyW6FMUwYaaQKd
+mIonq5B6JEBMgCJoiyZ4FyEtnPV/OiwC5mESoZQcoADuD9IxwC7s8LBDeKsq9L2NKUF8GHUSHNh
enQVssOPSZ5jaOZhvPiZexXKsHdxtGZ6VxK1La5RmZGOwQw/2GB30t/8+S5KFwc99xcXMGPc2JHl
39gYuULWYQG7ZEV929IGut/wKRwJMH7Py0QhXcSMxt1VBns05xsmUpLbBE5k05I8GOlPH0YEAHAo
QEsdZc0Ox1bpTujDkBrrLXnVicao0eH/NUg7Ih2Ke5aQvqiVPE4Fe1igO5XSH+IW2vAJPxjZ8aKq
Zhr+T3M5WNTA7MBoUBEivYikoe1uKNgMfbNsGOtmJ+84idxtx7XREtn4DtoZLYeBLYmmh39a469+
twxWYRCCmphpAUbTEIcPySFRzn/yOzkTpOTRr+XFz7/GNG3nBtEy3lE5u7olyyev1GpyiM7eQRT2
0tphCkkE5uo6fafQQBa9mednBxl0vmEbTnPQkXpt3xczFz5V1Ks/dOsAfktnNYnd282GhN67B/KX
gOlR67o4/wOxwWEwfhXOMrS/7HzujwV5eTKOUQDFpSS+WbpDVgmzsDmXpfNVRHDfLPFYqnh04D1Q
6NSLlVBBw3npbMxUPDc8Xy0mXKkZ0AoDg0LW8WRRMfuqvPzzgMgH5Wj/EYLFJkGtFiWXdjXiSK3E
iGr+ZcROK5fnwGtreAMj18FQoYZGJ/dkVMBFF2eJJbYEyOY6hBrLlBVJI2u7XO7sL/SVNr7FIOpV
87HxBTSxBJtmQvL1AUHb+am4M3ZgVnpfz4CQJyH4bCS7Nd+Ejz8EwSZlCa+g7s4FUE5w+TBoXksq
Q/geg0nT4jdkIcc+7Kt4E5eC+nZTw5riWm54v8SlnS2PnHGgZ9PFQ8klXdQtL7b/jbsAnPeItYQr
tQL0+fUBgB9llHFaTLQRrbTpc7ckVZF0xfzBm2YEBcn+4OnbhkciVImKfdCklLLaiX9ZbpMtGOll
BjAniybVYLK/XahnBNm5Kd99ECWqOCD7hartS0QMc1f2aq2zuN9CtQ553RPCrGouRz5sn+Xe8YiD
HuxZyln1CLJdYhaRMakuMgjUlEAer4ws++96qL60zKQrP0fS43lQlAGZ+zzjPtxWVczTRTRhjY8e
Rah5YU6qIS/8r63K9q+lpulHApPcxYFekzkAi3iM7tskBCCkglwcnVzYrz7zFjuHr63J1kSC4MAY
BkA+1gUPfJDBmL+NyWgcy9vHRabian8KeMqpzgPQMGMmwaKUyrGNG+h8a0Ny8vZZliWESErewhEP
FXYym9qQZ1/p6DKc0Jkn3Kxe2EwaTmAcvRxI+bzqqGCV49eybPlXDoqF7XztZtf/NJgEhaP1HhoV
Q899UGR6ipG9IW8mTLbUsyGD6wbANoj8WldNXI9CG+H02Lc7SWe717HAbymYWHawzAtEr2mPz7IQ
aGwjXBcbRA7H1447t7ix2AYCetLV7NzjF6zao6qOn1q/Im5F1uzNSn3BnKAGJD3FNeuYs4GEbQLZ
h6lAcAD9F+NMGuSCAVtacmXNc9Edn8dK5HOek3S+BUKJFXfcI3Am7E0/7sqJp/u7H1I60nFa2m5b
BMdraR9HT87MUM0wrrwkjHDwW0MQR2nYdUOzj5kJ8D5T9wOI80mPJ5q32dQRF9V2johLTd/v0KP8
zHLMYJbeAm8O2TluzrsdB45wyPXcmUe1OJLgWeg4InYhfWRHcFfSJH4tAoUpBFTGixQ/dnngL78C
39NSY/lmxb0cIKmu6EljO+MgKwtyW+x10cwQhvkuqmETKxALz9gKY7Bw6Fd4GRi0xgCPpFYrydeK
e7HV8Oe5S43bQicg4CFYeyRXac6feUROlh2A476z5ScHk25vpV/yUzZA8Rsz20/FPDxZlw9sfrOJ
/OFZ/HJNgVl++IjsYbldrZyM93TlZNAmFxs6zGbovsCP/8A6RA/i03Dr5gNnVXUO0+FxuUFgGLxy
uXvC9FyMeF7m5Vclj4fyRNsGuns5w0lljT1Lqb8EQo+u1Jx2gFRAiyzovxfl7yDbd2rXgQvmOP5A
C0wfQe3cBA+7xIyneDrhgBM5wqXefvmKmpsBuQe5eSC+4CNLxjrBvlhlzAYRN45e0eJe3pO9L5dQ
W7SHuN2/ZrT3fHG6YCUPv3+OSSt3ohhHzqCckh7pJY0wSRIhulK0se2BqS4J/+NWfzXTWZ9OjHrb
6Or2EZMS90Q5YuX+S8j2GF5qipCEOmBLs4cJV/t58V5vpPeh9w6nfpxY40M+Cm4h77EB73Nojx1M
vQ5NYBMYASd2GUxkUfXK3BQ8wUXK2uQrd8HRVZNi82RRXlng5L+N1cXBB1L/fg7Jo6/kGmHkOWrD
CwwF2mhlpnYuQPiMlcvU75bHl4eCL2sNOfnZcgBWyDU9Xnt2hfPJWSaATVKQ5zp0MwGfLbwvm6lc
H7sxf6Dqvz9K8bEyZfDAryp1cru/r0DFjfuViAOF1bVyor9eGTPh8nAgXmH5T/DpfGVeJ4sgLL2p
YqAfWnVQ5TpxUJCdX667bCpDnzVXnq4YLewZoifLL7YK0SIPRbCZTvGCpNGyu9nZqu0/vJiYGTXF
zWw+cWVsId2ORktBZ9KtxSpy9/cU8jF8bXPIRGPwHiDDpnqVHXfH4EQ668ATmPoDRXlKxJpSctYu
RAaynkCiyPP+4ZMyf0AHpe/7W1aSZ0a87vX5cAEZMpwk8OJlK+mGc5bKiP7zvGv+xO0PrObyWJ/E
IvHUD7U1ebciyz/B7ekT/eH4CwPP3mnQehVIzGaXl2u3cEmo1NJ3Lc+CUxUGR448XYMaDeRgwOSR
kE+BZzHMT2FtNQXODm5RnUJBIeLeEACPm61tZMRhqXPSSpIrKbiO80jZyDDjWDujCuOotA/kNnzb
VkKh/VpnNqnMDC+z5n5lmGc7EPJGPu+fJ3MuPvSiTIdceZmc1yYwh8zM298ON2p5kSRljxjviiCH
9LHNeOmqHIhdYoaQlpH/KROcLPvXv3ZhBQyNgrhEt9UwR9mxf/yHw0JCMgHKBAiKfwuYOKQoqTvz
bVVZCgaz/czwdQrneM9ZXRvTqWSgcrf47fXpc19VTpQa1Dx3gnbnqsnwinGBeEELJpppeN7WTfh/
yG4PNeVpW/uc0JECw2Vib+ALcE5nLmnSLCeTJe1N8Spn17/6wi6JMx5X1aZ3Et530CFwPrA99zWI
ftE1pnhJwzhfyP8Ww4Qta9ay22lm9l26x3jvGlTDexURw9+8TKaQKbflZV7BS0U2guXvQonsYUDl
QlhuqEHO5dXvOQ9UjYTA/SWsPnL5d2DV2Hj1ps2iW2l9tx+eozoi16mjaqXSMnOz+Z97B8NT1LpG
FrWfGK9pt6pd3n6biwBV2a3SAnZ/XUEe+lffvAPIjJozsScyd31YuvGrIaHGsvAFP8PkuiBB+UOl
Xu0U94U19IAKXJhblQ/dRlPZ4uIw6Y0TLAOE/01IKlA3Imvb9U00vBO3INffPZZung4UM2Nt8Mi9
srDYzN/joMX0o+eX7ATmT8nBRDMP6ntNlh1LfqgLDJAHwbMLIoCu7yql/CVQ0SSgEsGI3C399v3T
feH4/ZfQfPGKaXhQAoy2qdXD+tPt8stAn1t/Tto1wJHtTjwgdJjMiwFWBxaM+RSo+gMLzVYlAKH8
f0egPC3dntFx7rSftFd67Ubxsf41iAIkNVrdzWoK7NDV4PIOpvEab1ZmcRNBTIL4LFr2Q+Y4Rhbn
2LtlKYbAvf/Gc2NeihI9zPmmnGges+Dvc/lku6X05wASy4Vcr9mnOrFMby1kw559MjVbXYS8P16W
GgrdjOA1IUWyzFmY7ABWlxHB5n3m+HPNHJWcwEN26V/o2Cu3O08b6K5HDubn9Slr5bTGQKT4uZke
6iEeR6DHaNoeye2Ke58+goJYgUB4+BqZlR+YKhW0zL/ILC7fjIvG1O2OdB3j2VNkarHWvGnR3rFe
xbRFHDvaKB4yCADCXHs0jxx+DqxhmLYz+TnVaxMAHw5cx5Rgi7c73QXiGutsojTeuwwvuTpBcDDn
Pvpa8YGBaA9PUdYb+xIvVE680jX50jwaBkSRiHbgIY/QbElbvfmItiFmAwsWhjJiD8XpaD9f5Kuw
8uVuemPpmbfW4j7tbOqoJIKnL9M2cDbPk73PUFrU5r7RZO4aMa4gbDmtOkxE9oyTfQYG0kFYRP2b
GG4zZ2TlnckFnKrmuS8yYK+LyR9V3vsQztR/RUCeiAN11jdKwdBpePfMXwuYb3vvy84H+Wuir26b
5ceTiccljKIvvs4iaBTIwy7ItnkEXp/jb02BFSz92j2Sm6v1MdxQTBTdfEX7V4lfwBW4GylMRUf5
sxzrVDIbRkX2TT8AtqtEt7Irjk6hV63EssZK6KQyOaGgO40kSgF7sIxOCzhv3jH69pytgvaDsSvH
Nf64ZZKbFjVjaT5XLFmy5qLotO5wWra+siNZh7qwnw2YCjuCvjUfKBt5h3f2X2ifprMVTSiNdbXU
vfF+94a32OB2c1Y+f+MkwqjDOYfTuDiJl1PMS5xyesyXjz39lWA/f5vpK8ZWGA4vpWfYuUYZJ6B+
WzQIryOkZ9adVAYiIiSnSrFdXqtdqwF7FP+2H6HSVPOeQan6jny8ouwWNfXA7Ns9YVhlMO31EpOj
6zvPPgyvMuBWE4/PWk1VPKkXIFrCconGi4J0/ZYOPy7UAneywMLlK/j1bGJAOWbNBxsqoF0jcC9j
6oQ6GNbxLes7sCqLEGMMcYklk4vMvVqa4zNqHXLk+SZYBPknoRym4Ac+I9ReBpEO2d0y9GENxuWw
okvuR16mJCF9ng/276JU5kZ5hyfBGrkqIn4KBp/4W8c8vS/Y3ysUuEpyT+yqYjXg7M5YmTaqb4S9
tvbeumXVk8SeX65cemfa0fbXUrshDMz61i3L9oMeWqa6SkRC+GZfxVr/izmBWH39dsOHvLQaL9m6
1R+7UfXtpNqIH8JbZLc6hxGTV9eZuylPYO9vX8OrshyPihwqhCFaUcNAxUeYGCaLIBfdugee6rTz
Net1lCUbmHEFzfbGildWB+5rfIzfa05bBotyCEl4aZZv6Mm7He1otIs114hvcjCzqa5KBk1cns0m
vadjd4qx/XZqGCT50NKnceDCv8S97HVZu2mZk3vsjJJW4LFqp+OPWIQDd55qJ+s0KLBkZH5Tofrn
NT9eXqkzqXZQ0nfvfSOhKQ3H3Uq/taah55rNbuW9ner+50twfLBwRx6E6zR3GKTxyPiNzIe+f9AE
mr19vBOtmWXuBLk77S95Um+XqXam7SrakJyZOERbGp/3YcFFqFFXzx2j8L6NO5+x2kLJ4WXKpAB4
FgODR3q0w4pVivKR+FNFVz7PFmcom3Tv8NwMzt9NuyLiofuCsDMkSuiwmcEb3Y9fgLkC3HjyxvP9
H1Xs1K2DHFMrYUgGEZgd4GxFTWilKsOr5Ozkx3fiqZaP8+q3jynKxzxXDxT/W3ybat4E3xmvVrWS
9WRMWP/EJCNxwzxQDEHNosuKdlO9Vvwk0/dixV3ImwEcFanjsWjrCvBpAew7LuX9zLR4Mq1DSYbl
8yu4NztaJY7fk3rWB/ixY46pa9eII1M10Lrla4urz3Yv+N+Nkrdlqz6RF4qWgioJP9sPt5AE+ywR
82HkI4zeXVRk/aO14wGK43SX8q3RrDSGxEnfzdIGMhBYhA68IKcOJmNB3PspXtz7FQwAYyZw0ny2
TP8K7eIlNH6k45x4kR0jaD6gP3wDSF++ja0BjinGDJnlDiUUkht5BlH4QHclatFz64LvPXV3qZUj
dZ85ywjyOVDAhG/Gp2ebUL7ukgH5Nv1IuVeJ1g42HPuQFgvlS/xo1RUR75bWAd3WwdraWY4d1kLM
LOPkbL6L55xZjpNuX83z9we+JZ4/HzThrgfHTGJFIsZj4qS5QBFLUUFLpKiXVY/SLQI+H8QOYwRJ
tARwG8N9jembJBxx6kSuABUI98vttcjjGscTGirVEBwsCehvjjy9bR8XgM2SYJBEc4XsbeJ/ZqOu
TSZCtSWBv4LvKu1Hc+5IVSPIAKDIirveD344OfbRSktvXsCYtdDZgEqsWvER89T3/7MhJ4rRrvec
0hJXrXgTCHDMMCBnNfpprtPLPVJ6neMzng0V4wDRFu1POEVzFjmRTyyAiPuRNeMKq/wciy0QiNEo
asCg1szSFEBppr9SavwSzyFS0zsxqthxGtxv0dK7alW4d/EZWOaLSq4AEhwM1g+9swToSCuQ82qj
2VXj2k5XyCKnVt93ES0ixXeBxwtgiAUA51o1jSfZtONAhIk3b9MRAx6LVNL7lbAd1iO3Sq4ewGrG
aFiULQ7Kv9orf8sD22Ip/sUem12VZN7QDjQ4DWDKLTi7kiVg4u8h1hQ6J5yZrIu2vC1bAr27TcWd
FFNV6ZLkmEHJgOzQSI+SGiI5UANW4GqNahs2ok7G+rRDb2MvRO6cedLAZzFxrUyBpVvqN88Et+uZ
imuYIEv9QGEjrdGBdhGB1Pc9MVnFrBw07GTVO3IdbIgAoOuDqND6CzNTwR64yYBHY6EqRZToM+NO
reAMDVIhSNSh3sg3clSVuk+e4c0rqdiAutTVgpdg6c7BhST0zsuZYUwvFckQvsws8nlUqjKY595I
ZEg2XoKRG+vtKsxSxzmSA7kdrMjzAgExV/MPA/v8q+fmjMCAZfx8iy0kEmcLoCR8OxWU2ZU42G0K
bVlhMRfSi8RHVo8G/w/yNdUoT8j/Eqi6TXQe9m1JAqst7REzkwly8OLeULByAeHIbdekD6XyfZl5
3/aceeDOaPJTnmR9TC6JPw+7XbC+VaZzl4nVanGtkOn9fqwrwN3HLlatHxNmHGquoAeYvRs3u3K9
aly0KMVWFc7FGU8Zl2y7QkRt3a/hlqHYNsPA6hWRdJDivgro+ClD2UsnKkhub7bu9d6jcYJEnzuj
0Xn1wGjnHx7FQCoulfEKmOR+FdQozWsCGVzQAYXWTlnxHA2UoQCkANbO+Fu9Hg+iXdsNExU2bAya
lIALIDYE23RfZyUDO+gqO7QcM3h/+9yjFPB19mztW45xvHlIrNr/K/xlF1jFMvlayOt59WgG+mA9
mr9hd5U/P1hSqXGqKt0Fd2/g/7d9W0FsQXdOPY/ak4lVdiQ0riCyJrerd6Olp72CCXpENs+ftxIe
r+U6UhZzG5tplUeUZ2qmtxbI5Eu7s834Qag3wd0TMbCjnvxPlam1B0hj+IT2Nr/t3g4LoCDkN+jD
t/Syr6gumTLGVHg+s/767RYI+p2wRzYFUykHJ5jGPFW/FeOmryPE3kigZKGBlrV4D1KObtNriTyq
+bcWgNgaVSTXoflilpmx6MbeW3yP4QlDB6DjFuU4LaSNRz3AryldZtdPhuvQJdMa6lJsIN6hm/hh
Vnoo0VrOONK1GgSp6VuSXrJdsMw25aSvZYLFMEAGy/eU1jwH6l6qalIfXs8m692xqICZkZjSRzqZ
vx2xXWSy0TLFfGg6+jJQXppsREX2kvW/293E0syyV2KomAGlhq13j9Qpw6lK8JFagcg4V58awgzr
25E9o/MhJ/g/b8mYT9ikr/4nAaiJC3QFwY2P5TGe1Ibbdj6Tkcb/O3GcYoUD+lfxApTgdDJ2vaqV
vQt3DqUveNXt7k6oYxxWkIWfSBnV4CFlxYzZFaMY3SnNGFYfvDJyl9TDmZuwrBhOwVtXaziShEsG
Ir9HSLgd/YaUYVxTclkbVqQaJg3SsCmzalY7+2XWw6pKhmJ6dkxe9M6JIkj/zWHAxsVYtW4PlhkY
CuvtjwX7qUMgjcyGNujUcbisxWdbnCKRm0O9QIw0Ag2HCAg2To7D6kp3JwaCmyg7P3wFO0zKbmky
Pg+kPx6PJ6bTXQSXfK8q9wL46cIhRT8B6wMZfLyhJk2/I60mmHxL9BwePW6yIQElnJI0mtKIAPFI
7lwjkTE7q1iimwWc/N1tgceoKayTWGGlgh8mpe+mcE8Ef3q+opgY27ocEkzXeXQPkfyL0HvLqNZn
HN7eoMdgBHuxuOyY1SN1OplZDeiq72/mT50E/FiESBMkR2szl/siyx/CfyaSlsm4FHK7+WiihYfE
9DwgeYAThNBlFCmpXsZ4eIh5lIMxefx4EDvDVDfCe0dVe/70wen2NZmF8n/2F5dhsEzGxyExuWF+
8CNLrsDYZKrFEmrHd9zJmTH0CnjI0jHYKQikfHIAKHxtsUG4BYUZgV/SmFIxHv/3a398EuuRy7Ei
6teCZMufUYLKxDiyn4TvxXCyVtC68yMdLXcQTBM6/dDzknQYkjQwVl2W/Zg6YiU8fEw2q36BK5tE
2Bj3p6pl/AYRxcZs0sEoJ0TZrqlU9egxv0byVjEHsHDVMQ3/vxgnV6yX1t2EFGlM4fdBUGHeyTtr
Oc58Eq17dz9LATpW/UBbvQyHzFTh3ewSd+8skRlWkPBdFytkGKy4HEs5iWxncaMCSB9fw+pIBXvA
br9ekxhId8hTiYuQtyiVPjn/MRsXeIdD1Nr9BkoXChdgLk+0BwDGxhKsBXoWOHhsraP6elit1PBb
QQZzX4aQkBHx7eW9oUEl898kMoY5CGb+t/8YqY3QbKuQjwYxlscqESc5WXnccACTRpxqnT6ssGBp
6Hcso3Qri52xGKZewcjkkOO/KsNK7x2rnutFT/7jmzY+jlfmtT9nR8fSdzMi/SDlxbgD5rHwnOGb
7iP087+ACTuUackJX8KcI5RFUW+6UUEtwUxfm1az1Ss8bAArGvo19aMvME1db1vpWTIENE6AJ2CH
5JWpgEDSPDOIhrYd+VmGR0it6DxFhgQ5+8TJmiV7Wfb1OYBtECX/Z2HmW7cXLv8JrmMrWHUa3A/a
GsNYEXusbjRjKgNThjxeO9ydgSbtEToSaBMHIl4CcOVbYbbKM9exNUMZMomb4+Jv84jDU7/CFj7E
3Ldrpg+yTX+zVgW9lItaKrn2gpGsTIT4sGUoJ2QJJPQz0PlU2VG06YutowxAuwKisZExClbDO0/1
i0077oXo7XqBe6Ap4p+DvuHyIuuF+1UP2+P00bFVA/wWsSeTxaRNH4w/kzk5WmmxOXWSFq57+lJa
Y9ITxOyO3E1WMw0h7Kuun1Jr1fE+qIao15bXL4aQODki+E+tRW3PIBGhoUZkrU1Enkel1GcyCLTV
OvaCs3MkL7Ewi+Cy+/LXyGqXwwG4xtNDUeNNcbZJGAP4mSU6cvVXF2Uzrz0ku6kAqxvb63mm//0v
Z7Xm/DOiiLQMGz1v/iDZ8ll1Htkh0MhTEYrSPSSZqI4qmKTO8TCsLvoVtU7vpYHGSTDvmT5Oc3v1
qQPMoaFvAJvROOeXZ6MAFp4DHXPo/Yje6nV1Cab1oa84YIoTuz7ZjNtUsfLcew3OC8xvdsAnVmoh
mkLGplnPQ4/6SPewM8FFYomwBKTq0bf8YjGmHNqMjSOMTJ1aYkr+KnAB2+YTsTAOkTO66qUNcJtG
drlMCJ4Vbx3UEYPcQafu/3trTICxbAYuAK/1c/aVVrRJr2Rf3krh9UuZ9QuT/7tKoy+cE+10LEQe
7kZqitpeFlkq5MH6gysVrpekTb92f1HANzdzERlq6JuxIgAFA4Q5EbJGHz1GPPkiQGh7mTP1O3bv
k+sIN8o5MCj5eJtaMMdDMdMD3FsOcUaTDZRg/Q7wiiY9T6NoXX4/1U8A80KT23BbGKpsFZMQpl4T
ea3buhL9neX5L1/nhuCUVjieAoVYcWw68Stb1UjzOZjy4F6E8Nqbfmyde7EOR3JXzvBoez54A/aH
0N2QbdzZOvxp9BokG1L9TYHSEyAnMfYGIsj7KRAkM5lNRPsTV1qoKQZILDikDmW74lzvD2IlfpOh
ZoP0u4n/pES0BBN/YYxg7uxJjdWwBNXUr/z65PygonEgUDyKHfuewsFszaGUY8jMx1iUfvUvkiET
HpyXR9yyOvqLZUHYs7ypbu5wuiVVBcFyJCsIeIS+6RMu+VzsdD04j2s46FWmFtVIDxNZDN4qXNxB
7EzcZ7m4gtkWX/sq9zFlcjtGGZSczd/wiYnIS8m5KKRDmiKT0aVbMIzTb9Nxl99G1JvcSaH3VTGO
h+Nu2/2eUxDo/eA+Sy3qtff3SmcJWzajRh4cgKvEkIVP0WF6ncaESQl2HwyRDJceNJfFUzRC0clh
gAm+4ehpaaFnT+09jk3dfiN9y8rvvQxTrTcb5sepMhbloipgC1spU5eozcDshvCaNYKiR3mj+8Cd
TjhJ8lqw3/kohOmm72bLy9XO9rcZwPk3GZ2pT5i3gyXhjztL6L9UvprIILkVI/MmtOcLT6Sbh1Dg
2kzL4cFxgDTPm0X+dnQs0FY6TbtgWYwK5ZsMDSwslWDaO+BSBDoHttcTJG6s2oNJTCPdZ9UxccTk
H8GN7cSrIHB89m2D2Q+7ksuTgCRKlXJx1j7QJX6WDMpACKYR607L1pMaKKgbsudqWZp17Je3gidE
hvX/GFBPnJijDNqqz/+I4H6LykYcU/uJXmagEjYmPSFkcj9cV9WNZxkNcoEH1U3/yxzVtITvDVoc
5i8GNfS+ncz4e55se3OvkJlJs58GkbhjQBCRhm9zqnmJBhwZI+0LY92j6npcWQPDvo+/vjDkL0hj
V+DQbPY879GESBgoYvtyG4NyX1D8B1LdVsxPWmc56p2dYfWzOrQ8gtIuXNhXDYG6TIrsWd517Q/k
C2oHI//y+/kDNm5pBbH0nsZVJKvU2rwWqUMB5i/niCIeemk1za7c1UYgmweiQC3KbIjHrutYfdLX
uUXpDZMW13HkAsd0ryO81sjn+sL7Y34IT+K5ZgzrNitj2U+GZCFSyoMTKRGNfVVbR59URzhYBdFE
wku8w6E9NDDdJqxQy2T0yjhKee4ZZmdZ2/hoQMQgJdp/Vtf5KevP/JHnDMzCnYk1dFPGDP9fyFl3
JgbJvl5SfmYX3Cju1rDafqkiWoD/SHd6aRCGLzQ70PP2/WqZ5edQHMaXCOXpbXVT8IZ6iw0rSh4k
yJ2XkgJqSVx8xSR1m1Q5JPO/KDoZBzk9G2c1w6hApQzJHI12/fR8pHcqZIM7pTQ1ZTfASeDX1Xuk
kI5ldUHKkgfAoZAQqcnCnyUI/kTVSezZYOuIishqTLiyKGriFhXBEwNTzQdv2pEB5kOnLRTQDsrx
OAW8mVTql9JoBngWWnviLZHeioqOEUDouhqPABUySEATsOeurRf3bDfYf1uN1qQTn2eqG78BCQi/
cLFkaM51HOOE2urMAlIvHJxTR9sRODID3JwFO3IDXO6EeTB/2ZrHICXs+Mcz+BuGBlJveNvEnPYA
fXWK8V3GEqAvxkUdpHhLyjl7bolYBtucZGmdCW+vc/9gKWZ3Cgt+PU78fsVPjIAo8pVreJl9G88D
GCGNPxty+LS3FT6sJQnyxTAQbtIVnqgUMJQG3+xnoFWK034OdGWJ2a0Uo25G+RU8yRgzqdPvBvFm
4SQthaRF/CFpMFTX/i8eFJvj9C6xUGidzY3VTit/jxkFP5Wr6It44RhOYOmj/EtfpNMa9WSiB0Bo
ZqOr0G2lytfBcA6zJ1O10rbZ3u0U5pIZMd5y8JcF1Bzxp8/xyhHZP9hceHEWWs2/RQvnPG3/Z+Om
KQeAzeufduAhSIyNcKWewN2sWYl+vgfa4Zc7ZNXCbX5HVuSe9fbZPGSIFSU9VFx4LSnBC7Y0FBzK
hgeBJp5TzOnZnz/G3V4l1jyQ0bUt90IKeqdzlWU89Ae6cZYoB6gj/Ma3BQCNqM0cFXwWMTMM3U9d
By3HTo/sZ2gD4fseXuvx8QH2jszo5xBFskFDgd4vJ3NWz1PuRp9Pzlj44To94VS/rwzRSyaiXt8X
ZoOn8GvcfHBDGhD+JUNHEsTf+YgnCmr0fWN8NqA2SzIUOa+iFZHnyr9wc89OSGfsSUTmfw2LMIDB
xFtHmQmy4wLBub4xdweL5osXdOeOwagJtyneBn+I3lJnzLym68TAsDSqeOf1QEb7oEcGvcUillhR
GTYoGtiXpcxdCkb0+ZPHqhsuYRqjU/bw3TFTpQ1EZoeyHBIcp3VpkTHVMHxUiLrM0D6FKH++WBlF
BgsE0M375TI4ChHuwVeAaxOa9bsQQ0Ui7Z4RdQZQYuW5b9+Qx1SvUFLA8LJiXp7T5szvJMup9sWp
0lC1MCpzez3Wvi/JCXw6FxfD5kH1TKl1Dem17tSQNlCrUAB8cUSxuTVVJVnAz0za5dVY/HtksCpr
pYrskAtYQN8dBBBcc9ObGeu1aanUqkq5Ceat1eSTiSNoM16WCw4AQUzEsbIpJum696weEyZOX+je
YXmYOTRdoooLIfDpwA7i8QOghHizQ2kJrfCDRmnneifZzS6ixpbSBQ7Pn252kEVBvcIKpz7tVrro
ScII7F39M78Xp6hGPqVsVPv3+6p0StnjZH7QuhaXSU3eFdIOu588jzC6aA/CyCR6nIzBfZgHM1qA
xxWmRPWTLDASahWRRiZzwhzhhdMKJNXTAmRnadSzB+B19MaxqJZWADASfMFkIW1A/zRv5tFFbuZo
N4apjGkHfy9TnKRmG/vCQqy/zXgh+3VG1sPCb16vICki9rZAmoGxF7iM5YvUzJUbNfx5CcsQTQaI
2iZv0fluDvotlnWhxx08pc3cDYJHVKXgb2KJ1z04PKtWT3dAY3jY5Y2lbGwIEzXTORq7RY4mP9CI
J015d7XXPdHb8LMnLbeqdMQ60M9dPDThApNC2y6Iq8KJwlXbt+pDThSo2QdFv8H4MKjdeJVm83rC
nYH6Flso/ypkByer+nZgggwUTIvXjUZDoIz99FxBycEsTJ/WZXDqJa0lAagi6Dhqnt36ZlfFdFLB
2DzBM5HUNoxYv5n9wsJMepPte1H7iU0ZtN5QGS3lc8gv5aYQ4tG5xsrrqzQJUHxGt02kg6HCyHGm
9nIW034VAtR7OUVCnHkmPcsMHkyHH9RfZnUkyKceXa8dj5nUMmBasrQD9yCekndvcTA8qXeUbKyf
lUmhOVzp1zm3GVsjk/YRuTR6ndx+3bYwNhWKq3dPucqKUm0IXcWS62nZpp65nJ6QC3hMA3KV5NfC
6kEjzmf0uK7YAB/pbGi7mKeWzkJ8Qe6ZRzcKfXGXb5fj8CjTifVdvK35ZiQzJI4EnHwLz9hEzBM7
uwXfIpCP/sha9OO7I/01s2KhUMYgajbI2ic4Nnb41GImrVTuupI14Rtyb0Fzjrme0MDi9VFEtVm2
y21zZ56mnsNYoH9kmrgYxmyzXbnktdtaWDKBYG1TBckWz+vHE4/PX1gQIYvmxb/URCLO5skZ+aR5
706cXWb2Rw6lWmpi8yyiMC6l8YYokOIG/0VcERF5zJ6zc6zuGRbiin0EfbjQTVn5Ow1K9ws5349u
mHiCEtzLF0eXEEiEvF6+vVowX9eixegcyDyHAVUF70U/8fMv3y+ivRtr4bcwVtQHal4b7l2/0Dwa
dr34VDf5WKClOuJJPKIAKJjUmPyjt/s+esU9JAgmFyrNTDqHS/BIHUZ1gXK2/2pU/snKCJoSiXjM
BVdlOvmFKewa+SHy7uzMBliLbLfyMAugeDLqHVw1Vo3QMhhojZgyuQYBTlDMddTnm4XbLLmI2Wbd
6n6mRqJ3Zc1olmfhG88OjfSj40EcYLH56HPrgp39g3e6PWFM6GkNPmjnmhvJWRB7KZyJi3/VgmaE
jtH44ieMzrMnW0AlAqffFkQNUVP4rR3RWFGZTvBcYWzfcOLO2flfAM1il/5wv1mkg+tUDN9yIT75
TIHGSNce5yavr7U/d+JJhIbMBoGOlQM/UUwh2My7pkwI8YeQKRG3VsGMZL0S52a5+CQFt3zvKH1L
ClqOR6F5S0ofrarjgfDRUwvig+PDPrNE6m0KSY26/iPtzvaCQqKjaeJGIb5rfB38N7aNFTSnXYJx
tjuw3ZXDGtgj/t95QmHZ+E6MWuPDPaJpSWkAB+jG93+YV94X6IktIxB+N7CIQ/bgSFT1QGaWWTDf
pxtQbJgJxgzqgRnUhOd4GBccINUXNf+4U7csKfvgN/AwKeNWSq7ri5/3EJ3JfW0qfxudAxulKX/V
7uBjJWHb1p/Cr6JPPb696owEo7azHn8x6LY8Xu2t2rviRgx5mOxxmGl6vnPF2qmfPDJKpbO4oMV2
6nDP4lRYChN5KCpMl748969gqCh26eFXDeQkaOTdoKKgC+DEk7BgB/PmWx0s6MBHqGHm0Vs7KaE1
lS3vxetyPGYr1keEuCCAbP6CjbB1UzA/s7qXyLzy0qpDuY2g5QpXKBvXB1vCgGDdS1A+acqECUbw
J5Olo0VkvrZRS90uzWnOIhcMAiha8PfCZbJpibUa60H176FPgfML030CV4csRDMvqc+qH57CUlgl
RJPeVqlefWVmIw3xYy9eoiI+u/JNXeUQrgNByXT1xXpeEM7w2Cj9TioobvOIZ9Bmv0pI5wvXM+gX
soPkvEvgEgK8ht/z8SNWUAoT7vp9sN9YuJhCm+xbHEoMWeK/hS+w8Fq7Dz2IeUkRbggyLh8kE1UO
wEoDtvkCdSj8nvGPDePfDgUph542/XaDSJbDnpqFvD4B5Dz2Mjqjg/nu2qSqNL9cLPHqNMzV6FpC
59aiReAXw4S0Bk5L6WG1LpmiC+V527KBtfKdURpoqRzHOEtdHrLD1xwmOqcn03OiOwuwM/0+45qo
zu1z8hh68PM+hMO8CLuQfaSYrN0D/RT1qeh2KW5ngQyT2H1jdS1lQ+YDd8OCcFOfRyUYm2ztQpPe
lc7bjvUSOolQBnhN5Z2RiGugkLmCj3P7/gSC1uP+aRZaCdPRFMymLMyHyaV2Mdbm+ErsXERmox4J
jdp8GIC0SSgR1OT+mKsiIJknNu+cYtWL4rag+8tRZRDdLtd/sNcvQ4IMr3cSv7drB+CfGRUszmWw
DtT7e/V7LEagbR/MiiBnYS0+uFuLtzuyXe6cB5cV6KJz3MbB73zlYPOp2KRMqvBm90zeQzI5i33U
fLlo1dlS0jfK1gesmJ69nHZCegMmvbQNmCHm0V60Uo1Pg9lvlh90CSNFeTDcUCh95xj0yHuU21lu
fNZXPAC/wf9Xb8g8fjJKS8W4gckaG1wEUNm6KQu6SR/K2tGU8tYQWBjRyS/QL3yrO7OCIk+fo11w
M8n7mirTuzM89wSTcFHlYQi065CVmq+Ip2nCXnZlcgajNCUzXikfDJ3P7/pCJKuarMrZnlYPZPG3
snqosOZVaGXbSy3ZRCMk3Vu6fJBLmwvoSu34DO2VqNqZ7bYOg/7OAdxN/oKSh/03f8wYT40BV6Iq
1ymSQnbBbwwtNFhQ4j7n0qCiP8fa64EvKx1Q5xvDLxPqc1Eo0JypQULyGEy7XBXuFZP++7rmIKsr
yrZnLRo/Y226v5hxFV1K8PfyM+ibqMi08j2Tb7M95dJTDNrG2YaNOwCFzLEE2xALjhmdSM4fsQSf
65yoctds/PwSHEE0FASRoxKI2KSvuyTCyiY8ExzPkrWzJjguA/IOWhQYP25ZLMjb5djxUhYOjxWt
SR3TvJVzZyYJY/09/gCm9r8f2+1eSGbym4lF/Yh6ptBNGYeT0EGVYZKiRZpfKeoaqaa5yN8B+IMf
GsVlI/CNoF0X/JfnVRdirjFY6eCS7+FFBWnNoOip4rA8NueEVCOQUIo+Ydh9INOMh+t+5x6kQ0o4
7TUF20KFwCdCGtv9E7ynlH/+mrD8TlpDtvcEa2gvSDT3LcNjgOPr9Kp2yNqE+huT8EMIdPdUUBUR
fu62Vg8c5rHR2Tg6J1nf5JxQHQsz8xvk8nsmpVFjKsQ+GrTLVnET526gmQn9jMK6UkpJVPTh8E2E
c2MZTFcQ06EhCWE5LfkaHm5ZJcwYcEE9PjCviCYe7SRbg+HU6TKns5Wg6MuuNs5N0XzY1RtB40MZ
H/V6JymJ1X4sRG4YaQs4VwyNKkh+1cS3pwGUoJ1zffhUxputBDnU2QJ94O0/4SQsar6Px4SKcP09
QafH7wIciS4e4treuXoNXe820mYUrQK55sCgikLX4GBw9GNKiMC6oVr2PFKJLZZQ780hxLSsZ/5s
SV5xzM58Q9lbGCqSvfqUCro/tm0B4YJw2XzBPk9p4OUve5eFpc7kNKCOKdptiXZc3Rh9mDkyZj2D
BgTziCAU+BOZzVaWqzkHxbsstjLvdyCuD8dBGo9gqz/yyIk0SAKVJq1dbxLa8vq/zwcd7oUnQfpp
iB4fPwrIzo0YbLm5Jvav3a7HKhKWQz0xRyPIJeHNhF4GPxLpocaIKUn97i4j5ktxpgMAuvM4BXKw
n1fbUSnTEqgEKw/XzNE+QztsfIiqlgJdDwBpdeUEI5itzAlfuJms/oSphvE6v1+ok4KCOXwlsjNd
KibV75GyViS1u3ECWzuedQR+Ny9F/sCwd6dSSLzYgILIagrDNkmDuZXphbRwLVYPLyDuccbIKsWp
h1665dkiAMcgf3Abauglh3Lzfd5oZ0h8NZGzSAy31/wljQLtRFRGrPGzcah+jreI90eFZGbkhL1H
9jdILRquO0eqMCP1bQDX6vMYDBi47I57uAiDNYkGCW/t6v5LH3b6kBYGKsZ/nZS3eqh6hlS0VaFr
FLTMhIi0Mbh/5Rb9ZXxeUbRNAji9imjS2TYerAV8SSpdynnKO8ABupHeq0/duTZWioXV6Qr79vcb
r/JzCJ+iscQ8ZiJFrO6YtHV9nu99lg9Iu4Ki9w4TUBWjAOeHt+BkKS7osRwpDR0gaSW/geS7wIwH
4vRKs3kEbVopFK0BmmblIAiNkZdEfGST8kED+DWlR2Hyt40iDPP3rqrqqYqPLUhrjY/UHc1o4Xgf
NwRwmNwlyVkKN1iqsVoA6xoyOcbDUnIDSCIKVBlkMT0SUXriLGyWiVLmPEjC/1GU3pyNh3orbra+
B52CA/JoYGHeE5z7rprr6ETIfWubsoz1+VxS4JTc/Qva2wlGbjGGokQfdIgJKSjEzoSPp1s+oV+N
gdrYIbH87nJwbRiNkJFqS2WCrPdoGf9ng72K5CDFK2h2iiPBYi/xhvtwtDkUHvSY7kfIwsviTM+K
BBF/lOd3wa2YTFdEOBcklQekLzIB6iUbE8UiFoueFfqhqakADXrtGiZ81IGq13FMmNchaliY9oAU
W/XCtuX9dBuanHTtXKFCu3KCPrn34nu1Y3TcJFR4cCYj7ugchHmbkmYL+9wphh896Bpc4YiY9rRv
BgImWhGLNvwKEo3SfKIpm5x2lN6WSz6HO0OcMaYOWJb06mvha4lhK4ejGGMdqy62I3kcPHJhADMB
voRhYdgZcLxF0qnlTP1Z4Z76RJIvIuFwAp5xp1iGHC9AjToA9h5dps9Kvb9mY4fxmIkUoXSZIshh
y8+uIGoaETzTHNNAUuBIDtuQ2e9FuUXXYsJwUifWZCAN7CzQmADgIEXPpQAlt1MI4L2vsH02uGLV
ncfnrSwuQYgcQjA1NQ6v5aPZ+66oCnSN2ro83MgMzq3qXaedYF/DYkb6dyGjbNZzFkFmpiAYC4wd
uFUApdtGja0tm/HGqLgnNa5vyDjmZRIYdPFpnyevt/cp2tk5F6fm+9Xx7AGBc8voTxINd+z3E/mM
HVNwDMHQ/rRu2g/UOOzkKiOxy7U/F9WmE9HwFVk7J20N5+u0gHsNx3PWWO4b4QJNv7MZLp7FXCAM
qfrjdrTN3F2YerQITt8dlEIaIGNnwwd3asMbJ4YbsYU2iIL954/LBPLIP5exT/TehCmQUS0sDMvV
LO9zqF0elVT3wuJl7Bw7D+Iw+vrKxw3YUgLQPFPDyHli8qNphtnQSYhLy0PO1zRQ1VzPSR1ILOPw
cQnSqUsNFVPJ+UUBdWzc2n74+vWoCyJqaVfT+Xy6CX+T4F7IWkOXDiuRkRhb9pY0t0VGYfXriieP
9hmXQbBGGA0NmAwQlAsAjINtWe6RubWQvBFe0MhzLnPqpD4dJwNYFrep5qzAp4JdG63/9BjZnjz5
KHlG60dyXuHxhugAU+MHZmBqcChQZQ7GYRF7/fvXPzeZ9OfYjmTm5jn6tBVwaF641Usiso6798tD
uv3ZLbt/Jg11vB/grvZUQabp/HG3o8zcQUbQdMY5s1M3UAS1mbSa3HLNX4duyPmzdU89zzgGa7j6
iPRPCsur9JMj9Fk5mbxcN6R6gNFbYAcbbBbuZxrNYQaEg+5lnRlD4nL1bG3i7/m4wHL4d/y0j00W
7GvqIwekM+5fu7rwGegCtlLSYqYOrJgH6X8b3Sx2tcFNsrQBJ+mhmsXyOvIe4SNllWCVou1oD4JV
Nd4H2NaIiXnaQjujfAvyOQwTedh3tuFIwz82L0QS9fmj+cqrHcS0jb1g5PGykCwOYgUIuEP5jwcY
78jvw8ukTrqR9EPCNnelIPMwWZ9LXg9VB7/cr8bQniQaygyeTKQIFZK9jbNi3Pp+40MoFdztI7Nf
PXn8qAsTHJi29MW394Xa6EGrual2KAgElCaN6rUDoW0AKCO3bWvU2Wtq1CcBhHXI8u1CmqQcDfe+
/kJ5pHBGYzSg/BFENF9sriazoG+KqngRideHFZjSwDFoqvxpZcdlxBDYMMC8h4XUxi8jqBO/jJ3u
u66riBVhUFLVR7t+4tNyuvTE4U/LKY13w706DV69Beln6y8V1YOMFFDJJfOLfwTpFLzUXgHCWKAj
O6CxczIQJiHDE++nZvPPjHnWizC0LCMiIBuHtA/xkQ8Bte7+dUrb3kCrEJIt4Hdpntmacsk/sakM
TYf6De2QfHkLmY5lZKk5KsLjLwjzSxCesVvaFJm7EciF73u/9EcyNPdRVCyph1Ff9SYnvbbUdphH
c2ZzG45Jhk+0CpBdmoeUbjYV07phT5bNVZ3S/asrG4u8Jd4x+9TnpeEnKdsvAZJnOywZi4W2415N
mX+I9m31o7dxt8EWVR1cGbAxdrDg+OueRn2Dn3odJjPnhVH/QntRHbHRBrlofDlaMhgslA6duMJX
R/TIDYcZCQNgYqhhpoYn34zC46l58FnTaPBLsIjRtXrc4f4wLac03CngHAG3G4S+/XcUupLKPiPH
SGt2/hSt+ejq2d4Rmcvc0kzJs5eRc2vu0C8pPeEOoZrlwrPIactvVm8LLMpBlnFaPg8jNaWsn6Gj
9HQb2wTOdirRN5N8ONHbeYXcqszerXTDQSjZafSXB7rsF2vS7/x+8LpGQW7rE5k5oREQ3zJIRaX5
7yyO1cO32oRztkgF2OgVB30GEKJnbueH6s/vzbqJrrx7Lbtac2FEPQBAC4C2f8Q5ImmsHmzK062u
003WE46i67Xg42IA2SKjPdx2mp1yXOcRK7oz9UhqGgS9mZ14jxoOwQ0qWPybTvckPfMpC5plchXk
Mofx/YmuPN2Dt4DOoF3SE2F6ReqGcuCaGSxvVpFuOudEH8J8+unMm3RZBWm6GuDkG9RF5I2m7nPG
7vxoGTGMJMmeRopAKNfLF2eIshm9+XpzZ+CZhWLihrLydvVq6qf8bo+f50Bznp534U5MuX5UDjnB
MNUK7pUD+wLuO5yIdbYINxciMJJ44zVsVVBXBCn9sB76GpSh8u5zcF2K5gcTRB2seDxlPGx8jmeU
Eh5RIObFIn7ETn/3eyM9VLdDm8amkDS9027ipB32Ew04jRncCjNAdtY8InQ5IDYwRvVOs9mzXnPN
MOmKfH9776b1aihSYS8hY9GBXhqeWydFBQ9zgK7gD80kC03r+5RmYT4USEeELOq25oRsHCiN1bZx
r7A7qfOMBKCWo8mNeeapgCsQUvb2z4piuPHXQ5asyE+dK73LGZLThzKV+kXJ2lnfFwkXSZh8Ynhm
iKB5BuH0SpuL9DhBtvZ9SoPgmzQN556eOErGBWu6YbZW1FBbiKpjTNqNJOsp3sWncK4cAkjNFAZY
ay9Q3lTI/tUo87ZNbzU8+1KtBCvOF/e+XvmPL5d3tIS1XbN39NftaxVEfj5otdnRYqqeMVbk9jVv
ja6hObK9MSXfhy89pPxGfzAgvv1qYmIN0G6gAU6w4mmU2jTTVaqQfaaPXFcnusCYbQkiwTogkzid
5ielogaaKfgROiPlSYTxsi9TGdCOyNKlJrZTHCjUkih6w/aLxLApSo670D1l+fkDt1rEt1kXY3cG
KQQCJVqJ3/ab12M+yS2ZiYNCD+D01w2h3UEmBg8vtXEd7Bl7FezQOL8ZZs+ATft/4R+LDsk5Rd1q
amPb63lXJAWbsxouJ0LaSUAwmXIH4sLH8MoJVJJmF9L3Ky70gefwbc86htUwqrL8q0Lbw6uv+/CS
x69kcvRCx+JKnrnp2Aw6R9XnSKLjcx7vEGMMmkpb0cfWN4+d9DGr0cjE2lWPMTE/ByZVxgTKSCc9
c30AYLwRGruXcZd2oCbYSPODSwkkUC11VxF4uCPZlZB6HaquDuHhLWppGWGsPiblnWoieiKmAgQh
tiQqB/9LNuf/3jUtYaxF4c+HyB83VHF7YftbLx5sxBlCPVkXhPGcBLM2IkK5LEgLAwLBC6PRtkin
9s5wMQgAJW7aymuu+CCET7Tb/dWChrmALQCgL6blkupY/tuksUEfqvIRt7yjkOMtL4ytazV7D0Vr
Yz8pysUgsQucUJCcCyo24pKqjzgK8lqgwyDO1JR2gn8w88d4WygfYJMVEz2SMJWzTurXauNUT+E2
dB2gX3pv7FcACfyUS5kn2Bn4gfO+56LUHD1+3amSjPpYxHQMpfvQvrTnGbMr7hLW+Q0djX2uvOQ3
AnZkhbbgV0OmDUqKfNmk+9acEdURr5xn+qr3quMCeFaOGGf2e5CtxSSxTixREbTs+6UCnjhMDQBB
l5bj9PwxKor0rBI1sE+gqh460LE6o8KQw0ocys3MutN8LJTJvBHkv4z4ZgLmQkHwT9wkKFhEhVy9
H2ZYmLuFXSeS0yLMPSf+issbLeuk7nKJbUYBkVPVyXPd6jo9vMck77jXQo+DXGTQS4VqK9DRKDUH
buDDPr2bIPp29OUUjfKmJQKhsFz2llfly56Z5Am/NU4lRVy/fdKrN2GTqh7xuQvjKH0QwWxjqmss
LRkzpZuTiN44+j8UXc5/oiljwtzKOQ9osiQg8m39Y5OHRAKvL2Sy0sL+BsVwiAVRz4E6ALjWCppy
kjFOCNgY1yFF7aFr56IIz79kQoTIUXR4uQiWzzyMu6o1man2bQNt9YrfCWx+QscU4AlARDcr0uNd
Lwy7m5t/Pkv9nvzwIfwJKdQ3qQ40st8Rg2E0I8llxnb6YfBRB/rBGi4BmLlYIRVAwPCTfI3eezch
1VnjaVyEIJxphnJTKL+iHtvLLOEW5iOlQfZjFS9A2GHOZ0CV/21JDHUrrV00f4eFAx/8tSMlvx7e
6BqsvPO/6FA9Alh0yEy7VkrMVWnPVYZUif5mlDjHv/refVfeCAhyo/hEG9yczZLK8EJfjJcQ902c
2AB7GzC3BXs//bVwvqPDcAFR42o7/97CwUavxFDtl1JsmTFE2HE0wYWJx8nyzL1pbUcD/AZG6omf
NR5IrINEcPTXGSqyMYASpA/zR0/7jgKvRgWOG8ScPyp9ZhIFrhHeajKxQl1AyGN8BZpDUSis8NyL
NEDm5N0nFV0zGyWVLFC76eFTiXfPYHJPOlNL50lwr1CCW4SSqgjfGP/uJkMc3lmW2SqdMGkT4356
68Ce7xBq/pAFD987PM50BmDNlQyc7YdMjoF3T+cJkJxNWZuyhZZrtsLz1bKOhJaDcTuqBSe6AT8K
2XemPaAfrVwv246UEPcVVxG/B+0ZkS14rxG+LC4wiY79vk5zxYNNnLHZdn+A58+U8A9gfMWrhRYi
LwreSI11uAyyYxX/COfudfvCtnxZfGvCfDU4dN8jTeSugogshcPdfaW3xXSXUVq6DI+FANFP61de
Sn574iKupyHuSF3+/WgbKZGrltYlKbpW/y+K1U7hn4zOP9+R4AWq6TdEsVUbgcwhAa6pFNtom2VQ
tpMD6jwRTgfdnCpx0plVDFf2mZuq5H2gNssXnkPjvlTBQcQnyemeCt+wSrV6EAT5XuTwaRGoNqkO
w6nOpys3mxp80i/XeKhHjwlDZFA3WqaImfhFlr9tTlkkLHp8BJ6CWR8yHEsiq5WrdQVDIg2omrCl
OoYuSb7rBkPeNt8Xn9NiH1dBfL+SPoiR/qVdDn9htAbf5C18bzUeN29rTv08GcwPQXlKgsFzXtNB
K6tKJqvwcFnpitbzzeSGOKIhLxfllKaeDLt24qAGqe9dw8RdDF6mKdpEVRDF5KI+FdjAfQFuitMr
pmpFX45aUGOKdLp825UAAYjTRCl0syzVv37zsrMM+zLgN43tc4lby6TKBOe/cBuTFrtiR+susfaI
YwwpSj8Jed0LYuPz94KpX4+FYbgPmJRIGQv+M7OsVwyZIqO7nAbsWyprmOJJFXZ77zBqpizwzxqu
SJWuuExV8MQ9+c3mFPxU0+fvwqxTb1tD132MLJ5Ql3bso45BQmR9Oa3UwB/9wnhFE03rL+qyp/KK
OoiHy+dK6v5vxocYC+Ffhx+U7cvxYfbfSxxDz7eu75V8z8kDD+cieVZvfH5xWuyPONUBnJUkK+tQ
lU6CELYUsTcJFu+2pI7XIwyfMZQDO7ZPW7alPq3EyghnzYyRXcOsEQao2acaJ2Yq/APSFI+JXm0y
qApQJwgASEVE/gmVNnjAcHeufgE4kd/+iJIHy4Qm3mdGMMcNWDLrCFsTCi/7cpl/xMmaIjzE3fVG
rDhecWqnAiDTMeVWtgPCdikJAgf/OJ0zAADU04lAEJ+clxCQgOzv1Kc/ZpoHOGwPT/G4kwmwzjZc
o4ALkdCYMhr3CFeAqPLq/ht2Ac5TRhQVegxQ0A2nK7038/KJ8mo/VBQ+uzXwnM+B0SO3O0oaP+GS
9E3wx7WtUj3PJxnAj5GSiIRNI+7NDiUUoZPhy0fhmQqaEd3oiyt8weWaWyK63oYKGMXfET28guJ+
EeLrrhxx3dsSkYgsaJHgI9Kx0GhWi2AnouzkAz12fehrKXHN7iL32wJ4x0DtHaTMyb3S0IuyUuBE
p0So9JC6jBVsOotDDykhYFQZC7smuEulHjV7yWJFBZ95BZD4UdcMvpQZ6pVo6KfB+lwltbv7QMTU
T8/CZ6Z6G8Q5LSYXbr3sb0aptQnOP7FxUb7y0xxS18JPcm3zQG4NFNe8yPQuzhKWLn38VMyWgpI1
W2PRT4mIuoSTsvf3fESzlokNzkocVpuOz9YGOx33YSn5zWUpus/MRQxWPYl9BWs6Qsgx3Ri74d0y
b7Dme9r3jl/cxwr+DKPfd4DZ2n1tS8mm+5PlwSB4qH1GvRzPWNwnIBdbMkzG5x3QQAALUINULKUi
voskG3o/6vf8Kjb4DsMJt103jfNGFjxbuE2BOPzEBilJLBR+Lwyemq4eV/ZeNih/fUcMA0ZYLUCF
xwmLVD/YEH/gBhNTpkf+d98eC3RTS1BHO48ymUt9pIPpaPX1Yq2L0h2/JtLCkodkRyn7sW4dkHRJ
2h56gqdjCggGjb4LOxwuhaGsnBor/ah/Lz5gS+abysW14ISTqvDh5qrPRFm1JhO6sm3iZatMcS3V
GyRRShsIyqyp8aNwkc9aS6I0J9kwZI2sW6NsN5ckdeF/0MFUeQ8NAu9px3Qcxq3ZSA79W9zQxNSs
SOJ+rDXW74ckUa79FY+MdWDxkMUykYIAKIMdMGxm29q7re/3o+c+Gs519fDjg+4goJXoI24dW9yl
KmrZ2NyzogLvVCMvzjLXDoOCFrywBlBhr6wbWcfe1hkJrm1LJ+fQGxgMvtq6A0ShsbFi2DyhWKSP
KYfDD8FSqo3+jMatRILadUMb21Le4TADSr8q7ObWVVhCrU5DznfGo6pNpY7iZ+4q2pBZWmzyObRN
bw8E1zEfJTOc8jKi1AX6+B/RfkQl5zGvVfvEhCGtxrTc7F/uyOrVbbV/V2pCkNNBGdgf/tyEM3kp
BET0TVAC2GNNLBB4UGHhkyoAAPKr4rlhpqnj8FE3qZL2UIcvkOTmWedOtk1vivuRRJ4bH65tZk9Y
UCGyVNmSsjMXK4m75cSFTqGjM9rrWaDZIcs4ZoyQl0rlJwCgoKlOJjo14IcJlAKnrshzrXue5f/1
FzxNuFW6Nqqht2cK7I3y/7CVlsJKF5xsmIuMpbv7jVe1z8adJi4VnCIhoVLOfp2iXM02OoFNC8zT
zoiuvSgjpgsbFWVA1AVG0PBiJ0oFcbCgA0duuc75CzjBsGf/Htw8wOofNUfhL/BM2bcCseKuXkf6
ntHIy3QLKjII82t44AV0bXZM/GuvvaSf0YxmDi4480TaD0il/3bTcTo+SKFE/PoP3ZTB/jJ+vS5G
sLpcVTJh+6U/XVv94e2Rg+2AgRX7BdeH4r/xBonhfLnRmcUa2b8vcAYKJQxtEdjBdH4WFsMzQeC8
2wIlTxkpQe5QDaMRmyKmjYq8ihVcJelRser+EVqK6Vczbd38JihqSrixsUfqlAp8tv9s4yY3MHRg
xwIuMyyrYPRfCSEvjQDlbvrXFeOuf+JOSU+bWD40TaBDOL1hmCSiVJ+utrYwB0eBHSe/ws7RGamF
E+QVvukUzHjCvce6Pio7ZSmG8yNJWhJC51A/rzohkpMq9V2ZUSLxZMLWy6+nyY5iCUH40il3r3es
PG7dt7/OUsik1Iff9zlx0gXysO9w7VPY8KRnKLc7/tglGLcak42ZszXwG/EM+zaohfLbh0ct5GXl
Z7JwLynPZSwsMNZRNeXFqNrWjrJs0GK87qnw/2FB0GuwdSZ80ANrkOhBvhQ+H/LelWFGSC1OwxoF
4qtMyH8oDCKRRaI14EUbO8M5+wWOj1/WTbG4fnSs566Or/E+I3jNbyyCc2wc2oUJBVL6iNQ6SqdQ
FQOswjgG+lsah5K+0l1TpByIvvZ7rYy330bjrYgchUmjuMyMtdlMMg/ERPXq743IU+YwfKmdEtrp
7N+xfqGTK1F1xXscdWN+W27FtY5RDxLh5hvwyVEazo0icyF94aqcem1424ICyH26YvL4260b8cnv
1tFmYJuFTPCcVzQVlT38mPB7w/PIYAhWsm5t66YzlZhb1NDwMzPz/zmKqYZvsbIq8Ch8kuyV1Ejk
rTUHVtqkLth9zatHQHkFcQaW4y3zKpnmjbvqbvptKVovf1BGVedlnpymuJJgPr2kX1e/XRhpFLTX
q55wAohYMrYP05Tu9MKZQHSsVrJUIYzKZCYu/UYXppv9z/I1YT4w8tpfYzjCgWNmPfFrx3vwKEOB
+X4KM+/9602LRIopfPwd3qQEKbVtgZNeqJFf3XfU1IYbeTQnaAVELxYyQZShIJqyT9Xj75WGMiUJ
P8ryor0zoMh72mDmWP3nl/5e3J0FDIQM2M2unBlgQ7v0abvlmIUswDdgm0pTcBw1bxM2rg07vvnQ
txUzzn/TgjHxrrsvup5K5gRrRPvHGLJdK9yvu7cxpHklYH4Ak74OYVgwqyEplGmfKFlYo+wRqmhJ
ETDvTrrnA2lz2pfEhcAWoLiR0DLJ2G4uAdI0tojJNW6pHHRsMaL7gZfkqfGIoVdh78kzBSoJA2+E
5ztwY2Y+tZnTHhaT6WXbMTaNU5ix0NMfrj/NygCoDSeF6Y4u/ENbVmNVrsjADffRyMgLwcEdeQYv
GTbFHUZZga3q8G67yWrgrm4A79c96gawwI0G/v7dcB16lw8lfrpII/d77Yhbi2nm7KB1b3P+4Vo2
aZWB/hn/a8chLkF7aHbKN6wMHDil4I9ySn3EXH9J1KDDO/RsCSBzV27hG+zaorxX4X6QpJ0ONUeq
CKotzCB3tqbfVlHcpWLynerxW9BZQDgvowaigUr3b6QcYD7Xg4MhXTDaUALd4OTRdKglTqJtGeU4
u7rTY1lN7Y3NwR/2tQAVVFd+q4uJGt/At5hd6kOUJj07tObU1ygT8vkrNzLukkrrjKjUEfk7JS7P
3XfWbE5bgGl8bvWEIACsilVRlrPwW1P9ZXr9UKKVoJ8cLG4ylxKBAS5zMgo6oUabOifqp0IEAPpc
aa3ZZEvQu+3DCZKSkIIr7d3VqJpIBtj3puK3roqgRWDO1ehZG0vKC96nMvCyFYSKCwwKTC0HZtyI
iL4BdVxR5flwwrg6TM/EsDLmpJpMLiJG3rHxz/gVoL5ccY+3HblPvojsxitoGaTgDjPmW3f3FD/H
9q0v3uTn8NBPSPQil3VFowAlu7cduVwHD10l8hCpAk3ipSpQKb5Uz9Kw1Nb5XlBiR4EOs3h90hHe
fXH8pVe2g/1fWZc8ABNLsC0gaqLYaXn7eA8J3OErfC/HV35xc+r2t3KYHC7fw8tGqyzZwyJrawh6
UKnq8lPkaRo9wPLvB1fujblQoRklAN8yy+LfStSss5YEddZBwifvwIovjDv6gMerEflpk8DE5PtU
dPPSiERTmE4heBODQb9XnUzJgzlPac8gqlcSpEzipDM1LsRu3bb+3UiceX90uyIlxb/nfl35yuXv
1aFRb1D7FiRUc81c93gNLgiC+LCPnAY+Mxsxn93pQQ1ckAKoCta+ABDR83JR4mUrSulQ/AknEkuG
KFvgGgyVgJfUQjh07XbocG+qQmEg5hCK/wLqsSAUmm8iFH4j5jV2M//5I2WmARubI5XOp0v8kYKG
XQtdMbBRgazqcPd3A8veZUr7TBURA65Z3fbYTwjbfmLnuClAFIRt4zPY8X2NTJkI2NurwMToJ+AJ
JVV8kPyjtyGIBSOcb0p09lAXsAooX2z65Mtt3U5S9IPt8jMpUML6ewIs2AfShEwdPE28n+IzHVeU
xu1/PJNtVMdeucYOJYTa+OZjL6VCsvGsSTzy/K6/lcTEgRMlacwN9HapaCq2x0LRsLuZ3S86eN0T
H1R51SvQvLQ34gyHEMF/aoULVfR/q+FojecweXwy5NBwhDLBqDSXcenwx1rqlrgCxZR83/AQmr/p
BnsDExDovuHH8capOBzvOh0nwI1mtlMSGCDAR9dv9H/H4Qz1SztR+ZE2Y1S86ORVAtaUwQGPICs2
NrA8stbOf0BjGCJg99AX63Q3UPMzuBdc2r5uX/ijNT3urQB8E/8oPlcmumuO7UMgTf5A0SwBH4kw
UfzeExgTBmA2Y4k9PCcJt4gY9XDq/bgSwTF1b2XElXEPrlCXrSXH0T1roh3p3fyNTiQtsXzQ8IM7
N/0LW6WMDYBdt/U6OQLaGOi6K7Cx13sL6xBqG8Hx/OAnYGQqsFm0/ULoMWSf75eXNty0YmjfbYJ7
9TwkDPD5+VYlc8DtrprvpefxhWe0BdqDQGUm7XZTAx3M3IXPqCsHshOSfrAHUFD2+gyIzokeSTZ3
OD/bKkb4KH2dlWLi1QGVRw0NXPUV5k1VsS2hno6DnQxCKPQN++m+t1FP/H80sq6cx+DWKhcl3aRs
6DwHt4Ehvh8cP+WiMpeMIRqzFMk9al7xFQgK+79eZe6umgqJHFi6vn+HDwzCEaLRMVIO5R8Ne1uM
o6HXUeOueQssympWoEciohdGzE7QSSbhN/O8sJZ4mopAXyB85IrhBD7E+10j5mAHDxCtrgtK+Vgd
V2RN1GN6AYVRh31fqsUfepSnVwqMuBuMGibMzAgXuBsF4hd/tinHX4VhJqvo83Qu/FIPTQQ/wvz1
dR4ES21qeRG9wgW9iKXOQDsKg96pHnaKqRW2CAw1xDoV7jIHRBzl9eOsUSv3BUxnZkzEc/lA86dl
W0xTebHdx6OeIjk9o4W0yQz/aX9DsBe1lVGNudWCrK+5wNgxyFC26hqyK2Td2LpZ3L/7C+5YzA96
L7WrQxhsApsFm6r7kSke8lT8eMBaoJ9OfZXmqEWeNr6od8cXsFxNDwIci53KNvrg2yfWV8l77Odc
EaTtew3HM6ZjfeuVSXsIa4fGf7DaI/0pbXWRE+CDRwiy+CP15HQpTwXdxvHxEBzSFX49YepbMDnb
pzRUajCFqeGvpfNpbnoVoqxTgE7RYlvy/mvdRE/QqVJ5l/mMdYrKLtt2lBWHkAe69W32ExcffuJ9
z9x3pK03rtBPUQbQXZCiu9Ll5C2xfAvTdFc0sFZ8Rqjxwf4NCxS/NdOXnVbR0ZXrBYMxU1VjfTnT
aMsw8iHMkbIMs8hP71aE6tnsGvzVwfxQ/LJKHWNxtHakW/RjP7v6Uwj5sT9dBBXbj5AG8CNoOITM
C+VWwzF9eXSZkEeGoyAivSnXBl7l4waHVrstNFNg7xUSnsO4J8KktwmXfUlDEcF9EapRX06W9REN
mE/SfyaHg6JiEJ6ByJsE1Pb1yBBE/7oZUqgJsickIXoFnn055mB7pGRFYvu37rS0iEyn5uUTdNHk
D37nBEi+tzfVTSyMZ/O3IVQUVT4VkUV/y+XHqgSRJxnzFqDAHqN9QAmhRhn2QTzlD3yqbxxDts3O
8o8KVOKMpLATn7GLu2Aspob9+l4/YFjDT4iixOJ1wxekPaO93ajU3qPyde5Mcr1S1fOFYnMCZ8HZ
wL+l/s13t0MKwd+wWsuvPGeTr5NgsVD5K0GNcAO/5uvBgqI0ySIVSKnyqrp1eHTSIxcNpWP3svox
P2xjsWoe6BQ2SXDo2KMZyNJxUm6oCJgxYIC3zT1nDQ+3RwVxTZbRH++CxWI7oDeuKCPDLe57aeUG
CsjE0WaGjzMpFcV77n5F+/JFODdrKiP8NPz6LkIMPXhIOGOxUtjq6ibBZncz6bEqO3O/O9x+jNE/
m8SmgM1m59WoaCdZ3DqtiH88BXV1bQ+wLpq5OQ5O5jIQ7u5Xy/Gq5/PDwiw5GW5soFV4akVC5f4n
o37PqgmQpiOGfyd+GzKNqk44QYTA562Emb2OhRPK4C2r5vlUagYkSw6H3YeIaBAznYMXeEwodxV8
jDb+8r7fiy8EvghZQkAmzmK8KmTBNHyWS292Bw5e2/jC2iMV2sG3wjbMFvP9dSnkSbEK63K332Nq
2knN4yV8xM/bvOu8rejz8SJDwr4xu24+0U+1zbKctktAL14U9YiA0P/qUmsyD4s9QpNhbLyr6S9r
7kvy3R2XRJrNnb2/cG6ewlNhgZsAjq2KNwxG/6eBrk3LFjn49Qn/ZCi5Az8bGPTiA8AjlCLy0ck6
6LTsDtZ60Sb3Nwd2rVM5AIUWQ4AUXkJFpYedlGgOTbhF2WHxYe8o+H6gq6HmRs4NZdoNJwSyywuX
D2XUzUqQ4OT2fzR/eCPmFJLQFNgdpIztsQNixLTyZ8rn7icBpqKXXW/NkkkB+HgVIwae6MpRw0jc
2jpD9xcpI5He17M8NMQQ+wAO1izG0G4zoD4XTrlwQfY69NuDMk1fQwixe1elm7/248+34yBoVXOt
yMbtOgatazdbb/L89q2Xtiz2OsTTZc9wHhV438oDewc15nO23F4ilKxobnK+psXJUUTxUDV1jz8O
u5Wu86TVx32xQXMd3j7t5BCrC0jO0XjaZ+xFsEpeq9C9MoKGrAo+a8uoWYjvG9oCZC7TvQ/6k6WF
zssyFblONEFH3mQKKUWrEJyyZnHp11KlLbc8e8mTRH7l64qy1BKb3SGIK76KEt+F6Kb7N8tyeC4v
f8AWRU6wYA2BvXF8MBX1eaiehbhaCxuJJC3/4ScOJN7GwtcQLJGPZ+7bR7Rr2Zo/iWHOx1THwi/U
gX6jn18rjmAWa8rJ3Wxj515McL/FDU453Tq3mb0VnCPapv1fBsIPOViRgMfBBZU+4Emus+jmDYak
VwbvP4RDSo7sjL9ExSRMnHiHEiYYSIBf+Lb8hZH6V6HnyEPsCapUBVelRUVOHj6asx2kenkQcZ6T
OvisDSriErI999YSQgY846iPzAVa3voCIR/tdGWhnkzMG6UTWAzW/sliGq5AccHwKJ6fqXRbGC2S
o8TnuSqvFpt/REgzmvkd+mlwHTb6o4kF6VWL83O4wxePB2WHPU6Isj05iEIK2odhW3gJPE2pf/5L
Z/cDYOCsVwncvjO9jL08c4DEhNJYhuJEcTXWfMObOFu+Kp5fpOdkRP8imnQeTwMGaAdgyETB+8dq
u89Ow8Z9HOU4MxogemrvC4BpCTaeavCqdS6y6Rt6NS8+2JmXNhpuI/PLNQthOhie+dbhYs/iFx1r
AzQ+sid7TixkYhXht6fbjNDFWptmfhb7X83YwjUgiN7buyjatQvHm5loSepic5kNPc6/l3bgMliy
c0lW7TciWh3BpSYAtZ4V79gvWh4N0ZsCch3C+lC5MwIImGh4iAfZ8arNce3QcVwqnX0RTS4rNKNO
V8TjmY5ntAJu8xkc1rNdMQoWumDsNH6cYw6OA+DFXnnwUay5Y2amdbScpbIs84KFXFTjO4bWWyQM
OI/FQeGkX/V4nW+U+5n9Ggwqdrfsr8w+VpS1FsA+h2fxhxAsJxEv7OfZb2qJqxsaGWhdmV7y3WcI
J+U1rKeZmtBcsFGvRSuLCGuFsOVGvDRIL6N1vZGvAs8Znc3PD5kFn0MyuN25o4I6JTX3WM/+Wg1R
klSwNxqdyQgFEoqbeN5KhqRljlOYMBki/xIv0a3BWWbi3JuL1dp4k+kLVe/PsVbI1m1yMWlWYdtK
yjF2ooLvhB/8UMCTL4rlzFEtePIpinF4RuDHd8tBTFifQuaP+cDQ8mjhksrHXDRgk5O4GoVw6ccu
XuxClbw7ohxnRSxKKcxrvGSe1J+6s98zEBDEq+pAqiPm4g2x6oxh280tNT+RVFedn0MjLAkIlTDF
l8aZ5eLuzve83Fidg8utiysFGFCMDsA0as9kzjn/lWyn9ztvHKtwxPu8876QIczbQGfYe4Uj0Cq2
EcIxaP9m4NUXOVFhb51sTf7j6mc9JzSFvQzX9WT1GtkbqSwR3/A0EfQPe2c+lo9mf2xUff0oIS5c
Z8Q56vfhGvhQCsviQT9iBxdMqaAS2+FNIfuDtkbM+1sl/wSqGhBoLpg7xcQhd3JkpxMg3g9uWtNp
Vi7qcDP4NgnSlvhA8aNgmZPESqblaOOPNziMTAD3qn6LEbfM8OhZ/LACdlWMjql9Ug4VOuh8mOBG
YnKWhnBWan2QZ49bPpowSIL5TwLViggbZ6u3GqHpP8QqfUPaNS5BgpGqus9fWDMFyPqOBtIrhUnO
fkkrkSb8CweAIpWHAmipFx2CJ6KnS1yqdm3gguks3PU/fwpztVDNToAshEuqEKWAlDv4A7gY1cwV
U3OLf1GQL8E0v+Q7AKdJ1FpW5wPj1vXSWo67BbjsjXAtfgh8bZf3hqmi3KkTTwCYmBT+PBPimIiv
L1G9gaPehDYTTcqnLa65LfaolKsAeeOcNOBXJmIdXU+yfwKRlPJmWF9pLk3sTp62WqC5FTgHVbKR
KUfQWHKnm59W+BDQeVZSPxc1x+zdHjQGtSI79USqzJ6PNZeDfVXu2tosc3QAbjR+3MxSHhI+dXQt
AO6KwzdE28jWRkgJTA39eZefMiL5beV7Up8TY39xDR9SvN2tbzi0IkONI4nwleWzboQtlLi7CLnb
m3+QCA5fUVi8KvzGtiGj1W+A0mXOOEe98nIFMFxtowf81pxTAVTn4KJOsur/xBuWFgX292vd9h5k
TuKYAVp/xliBdiCSjj7PGqPsM2FTFLvnMG09m2HBYIRCDAkjVSC4Ks23JlEQQsnZaNjWWq32/BUD
4A6Ly3WnlUK5UGu/7yNLNp2YcqDYjHBKF4DGmjA5BZF1oZNWA42UGe0/9VXrh2EJOh28ovHhwmf5
AUKsWYIkCemdT9sLyWLXAvPnZa9YlCuAngL08VSK0LiEuytNSxAGzlOGB2xxZtNDGJA5NfGaxga2
uKIx5OI1J7hbeQ5f2WZQ9cxZS0RPrTDQd+mApuDhUAlnKfRQDd1McNzChoUGZJ872H6tcoCvH8Lp
mG0FWuApaom6XBYsJ0HAUBZuZPwVqq1+pWEVF6JoBRScPXOaQYH+BSuWCol+rE8hwcWe78eF+CLh
jMZAEMcQ/vhe0VbLDPbLOeOhr+oK6GW8aBeimTDanpkJlUOY+ec5Ik/DHNZ01ZPqkK6oz8KWqDLM
ppikW+tZY6XPOIkcVRRYI6DppPEwGk3UazJTMEdSUE98+Xahw0EUUcO5/d/AclQObJLP9aG3fwxB
RKrqE1X4MJSimpzHF50lMkBanUny51kUjTnkD2CIzCW/i0P4OxMStf9fB2Zl30X1QULf3ymGx3UN
ULkwjJluab8GbKkbjpwncDkgzhQ5Ng6jJBbKhJt+kvd8quSaGzWZpyfPxDGpZSxr6B0siAbDVDpj
PDZe8bxuu0CUiZ0vCmzQqD9cELl6MnCyDLfWv7ZPLmzlutQfNhq8rhyLqHIuKhBxfMykQfSHjmLX
NMoziFA6cbh/UFNZCznIsH8m4ZnXVmt0Ltvj5q9huLZ+8egHfQilxnivffTmfve3H804IFzDJnte
wlPOgm6ZLxfeAfFiRhi0lHZU5btGNsblv9yqZcnBV+5cCGO/LqqsxPvlCEB9l4fbmpbomuP+spw3
JUzvuik+0I+NP8SdKlViiI/qeqg6NxoU/awH6gImzw+LlWo6oc/YCwl8Rbxg06mUaSkcnaKDoyXS
SqwlxFuXJKlbhdaFxdIe5gIOO6Ih56gYyMEwwy6800l0awa8fkEdBd5iQ1Wxt8R3/Q31nKUnrDXO
hHmKkx//kKQdjzOkJ6Ys8VAp6t9OKHkah4HCI3rPh6noVppNWcwwCz+/Hg7pjx2HDsOM7QpX/2qe
SpLLwDjELz7Q+eXW5QdN/tr4EQQm7g1ckthk/PpA3hkay447FOcuGl6sOdi6PF0l+dxFGy812zTv
62pqbzMZjyEzsRam0r9rzsqmeMSyPvhGQhkJIgejsLt7qAx6nyhJtuuo7reXPHonT948a1aLV4pA
lyq9mIQDPBvO71FKaVRsl/RQjxO4U5rhQ9puCdJr9V2/4s+TsXwIiOJl3ymbvQI9LXzQy9hN4wEJ
pna85/vS5EsX5eu+rgn5V4CPPygJFbMtBcbD6qKo0rTepIMrRkNVgXMQUwTjHM/rwJZJLtiOHZo5
MLqcs0VdOlOWggpTGLEnNCXiDqPE0Y4DNNfhkTt+e72Ny1k+PZLbsE5cOkS24usE9wDHjMj0PuxA
bIRV+8wnQgeE9rz0z+4/Xm6p5msD661cy79a+4zJrI+9NSgHDdDbWb0kVz5SE3wOMX2msmdfWyNz
nqfiVkHBNS9fSyZgjMSRRPW0E0V6r4b3DTOwqQ6Je+zJxcwDoinHIGOHsZZQVJUtL2m+eDS2GMG3
fybnaWvCOsIEx716zvwfu3qNYDLLscCB1R2Rf6yD+YRAsgSgSr4f0vTCUPLj5YPwkR1RDVS0T4js
5iJhkzKMl2J8ngq5i9Oank+xsXyvPjWab4XTrDneQbpFDNSQlBh9pLneuAu5/+3idmMwBeBuxodx
Lf9ynsPX5Hd83+Cy+qtov1qRP2uo6Ka6Ohj1cdc6Yk9LPR04AWN8pm4J5BIum/0UULMupD/M9Zc/
YdWBUUlVFai4XsLZ7BEHSb1ayzMd5e7UXhWoD5wqWPwBTMkwdP6JlCfRs8JHkwivEO0nEQ4LRrJc
AO478Hm76CH7G1Ydahwjorxn70vsbUNlqV3n9sku19HIlfeENATQGsXI64AiMX2qyDILMA3xaHh0
Sfulzho8+D+64MPjPbKfnuwMLO68UZbb01uwIWNvXI6UEZGV8ThBKM/3R25pQ2kzXgTxqIzGBcDR
b9wPedfcW84g6ysrp87rf7Ct6fpOl1WKeeB3dKRk/kn9/278SsLnUFsbCcWQiziPf3f53oL+O9e1
/BlgD3Dh2Cln4JIQoQj5Ug9DxhIPNOVOPllrKvw7sGctszDgsS1SFxAsKnoo2A59/R8pyiJ7hNat
01UPoVKkXiooOeEQ/ar7s452HDn9p9nxEASjIuvlObyf4a8aWwBR/8ej4mWvVpFD1uU4ohPtmGrx
akHvOGZvPZFUuY3dYlwiNGW8RvyB4fqzDs0OyTyX5FLHKpI5qWuwWvu8/wcvJ09blmIUrYCQNElw
I43WEQ618Z3KBDuKyv/T0qApmmfJtXSUNATgzALoWM8u9BSynj+hxD+2o7q+vrs/+ixuvj4+KdD1
rSnBgPMG4RcwlWtY6taDz9qWe4sDrNerXUXnRSOaqSzuaTKtC6wHdgY2yEnPRBHoLpbAX3WSXw7O
J51kzDq82vWl0OunH+r6q0LXUOM7YUIcoJC4HK1OAUfRyhfNBzPpTaiZqWyAOZQeHWCaFWXQWgBu
0unVoz7MJyXiMwW9ApVJG7bJbcV1zam+mjdbrqVr/F3HSGKGS3D01yLheIoXBH9uYqGGRmLPKAWw
vGiwlERmLLFZLXCjYWGVPGtlb2gNxQsmUDPMBGZKMeI0BEcETtiZlK/1s/lsRruarbMqPYa376iJ
A3OC4kRrsSEuaN3SqpR2Y5ryA4AtM3ad8dUKkRxNfoiqI5pWbJVRRZ34rCn65oLjbHbuizidDlDz
7U1usHY9NcLz0rhKGLUX23Zk4OCeSmdgPsdTtjI96pZE1vaNFII0tvgF0VzuKmWNHfCHGC7vW1k9
SELStWOU9AGPrpdqFxSEJ+CiM2IDCFrAj+Xd4IgDx1VAWhSY7kpmML+hesHZjHQqUQXSMPhEzO+4
PdsqUA6Q8HOHCz2TdZO4Px3iEa0S/iIKgRrkHFyOoYZ3Ong90OpRWov+ZaZdVbqQ43YqYIxy0M7C
WBLB5KA+3a0rgAs3vVZRZ/7d4LhV9pXuN3qNyXTOt1ITw00fMFwQLslybzmOmFJ9ywQ/3AXHbJ0h
9ySI/fd3mvzqDdIJmyvlDy4tI5qY/lNH5d1TeOa+ATqPniTapPaA9khNG+2zJxiESkVDcpic9nSp
WfW0DN2MM5+V5bxZWi5cWmSfuOh8foQQVBvA/I4TDAOfoiYBamvU2/eFeRp2FTLzqw0vCuOq40hQ
y1fFCfkDNEFZr3ieKlo308PDz70k3M0FTHBv9a2CMjPL59epfjmSgTUVj+bFoY911SL5yzvPlzXk
WxPnhIRB5RGCY2KifmGfM4QpsW9loFnqLAB+Dy8XyHYb7qmTd3djZQOBMlGyf5M+ITUnxO73dSBt
SqPXJYTCPBB9DTNZjMMoLTUm1j0pgMo87o5rL+cAqxRYiAD/MfVg9F0OI0DdJQsm34qRcy0FkuQA
8oyBIXzwicV30dVYoFGz3MyO5CGNxb/5iKZUuy8B2d94dYfJjH8W4meKGhrZUoIckjIuZ9RwT809
YolJcBgazNECe/h7SKyYoBb2oM5WokUWW0GrhJLV5ut/XVCANwkKiUpipqk5Ah/Ag+8X2ieh1STp
rCTsMvvNO5Q/ApAJDv75+xoPt55BOLjJD2nnby/Riercdy8UsO35tcpnvvCEke0EpBtZQnUJg4vH
W7gwJP1FjDhYra8vprLo2Z/pldnDJ8YZKXY55s1Jfx+PaQmxEDVQ6Z8v6aR/ttKKYj8FbnxoELQ9
evzba1ZmKt/uL93Z2Ar8sQ6/N1f2UtgVbTBnGrY9QB/pAJeDceH+9Y2IzpXUwUThtcvR0RnFRVtf
oasMQMFHjZ06QM940O4RSW3Vju6gF14qh6Z1ioAk3L3vytG9lE+8Dj4HHI6hIzPrt/Q/fHPAtjkW
lXkLYPWlmgIkJqgcJsJBGvJo3y/za45jMeWdhuhJQE5NNfRT8DqZ+4NwcopDp5X+brCO1G6r+phk
fsV6apMe2eMA4QbnoM9Qs0oWYfkHa+GypVqnduF7wNnOpnfRleGcW1kWF4FGhO6Pk41RdV8s5cIq
8HXK+xw7WI9rBxmnaC3Tx7Err1WCWQUWyge32O1ZOw1CZvtFIAqdnAGolZq+RgPWvR/VAiwF+Lvg
2bTAsaQ6/oIVxSJ3Y+MR5j8mvVCkyLxnDwrm0fZePhR4sIhLzcp5PlsyVS3YLF3zdeiEDnshJGZt
iRVBqhJGM5GdFcAhOTdFwqsAmnWMPDVb23oEivADR/jfnDG0UpLhnJ17hasTa2dsHwL3aw/0Uoz6
m5BDR2r000A/xVDjo8oyq7pM6DHRlZsDMOx6VVM6dCTnvI5xYdcnCB0/F4QEna1JNB/DZUIZ3dAd
JI/kicbeAKuPvfHhoCfG0TnZqf26SzXilQUIU2ZqEJgBTWBnCQHYFYrB72cGkYOQZrriJ36NQMdw
52LrIqGs4mGRWHGO51z5LNJawlNYUgJf9l7It6uzFf5r7w6qRUOLL9QBfLXgAHKx83+nWP91RHgJ
1EveunEZisT75fZnElSkWMO4iilkA12Wn9EmyaBEL58/9zwXDQOdztaksH8wDxAy/dclYRbmVrtl
fsWPTBUearySMAiDiHdDAuBBDIMfTLIEUynhsojtV0aXVebUETMnyfwMU80IAEUBA+HOhD7oUwgm
hUi8r9VzVvcTsc3jpJ2Da1CP1YEN+PJSpb90QwT7OLRU2D9IL9MpwV/8QAmV3GuyS0BWYvXQeSfs
/uqoJuX0JGCkNC5vPwmEZLsc14fAJ7mPEyFgdp05VCZ/dauhjF1poO1sMg/QrO1yLI88W9IiFTtr
ZttpWo89Rj6uPTgwBfTtQsVT/wME4ETK04adcf5bjfq/SJRZnEVtVVVcX9L3R9e2Jngm0/srUOP6
VXwNW0qz7oa7NY6/a8CPu6a16TcXHzN85TJnGagbsd09CkituchW+ySEBRXbTOr1kEP8B7PMlkUe
vVYerA+7nb5ywuGdzNfBYXAGT7OBIfBqp+Pr0+Lowr4UN5zLVvxc5cjq/8i64c0+z0cp/Cr1hrpL
H/YlBppmn74C9uzLyH/CZrZieSTlQnkn2CUctTbgzV5ZHjcT5I7MvA/XYH7mR6CrKphJ9FgST2Ln
HHxSJRud8J/4Xt+mr8AOq37g/ai/x/AkJLbFkg5TFh+SV2c8+XYG9ED5AzZGHMFzmHH4uN3o0mj/
7cSJH0Px+rq+dMQMd7nnQe70hsrZG/9F44Sd0AG533STXihXYLS5xHPkSuLVL3/gSXUL5k3T3/dr
z+tZjzTXsszM8Q32i0D3xZSLuTupvDLJ9XQlLBDTt7C3cLasUW7C+Ofm3ScAMk/7AyUC28+0r55I
lWhA/i65nwkjUOHGLG70B60Trm+sg6EsLhVuaIXV5UaS6UXTFQqsmXguL7nlcIpzTrSueAuwEWzU
KBdHIO/Aq4HtXPZJrRBbRwhLR7zpMOh1AF+Ei4FCrvQdJHz6HKLmqmN4QzrQwcOeqY5+jNYAiRe4
BOB0MUKEnPWKqIMVm4dvB7+58fujOEJEl8XNFsiMZmP2s4TCMPNMR/PvFKFchRPVBaFHkBZmGn9K
Nx9DhWcgzyse2CYt/WH4EheWm5brooyO5lbiyspXaEeFaYqCVv9ao1zPYVTlqYVkDE+VcXWVdOfp
8xT7c430bO2NGKNDSTeibyVLz4GFVVr2xgCWKIq4h7RWaGJeG+vsZd/GLhy66cx1GCAGENACaBwJ
WLg52kFwIdvJpSfaBgOZctabupKuUAyoOkZIVyBEM8R/kdYSKQsMJPfBilnwyrmgPvlkGb/Pn/n2
wGdifrJBeTAaZXbqrAykQK1kdfiNzCLJrkmNxsBpOrdecmd9s/eYbvFTwEuOgppWeE/nRLmtNPf9
Oo6TCb6shfsGU6C8DxCChm6RPZFUmd3/nTaeCgs7kN7pGmYvy1glF5/StUzCatw3gWF5ZOpaiUst
4xnZSRVN4Ifvg6ysunRhaB2TBCBOrk7lhchM/G8PsagfTwGAyclrtEM6Nd9X87gYSBjob+7bauVa
DRHa1YOa75tbkDFP84/iiRVy5v6wqilBfpDECNzUAh8/XowjOTPJ9xhg8LQWAbf3qIDAt03xqLrp
lx/YDNgdbS5OWBNfVOwZY1wWVXiDJSkbG1G4qov498nHPqk8aUsvue1qOHLX7mcpNqVO0q25r2I7
0gze05UxOgMJtqrxkDrdutoFeCjM445LhYr8hUMNVuFNcWPliX9Br3LKDN/0jJPYKR/T9mm6mNla
sbYXkWknE9bzF0M+tAbazI2JY3p0A/C72nnzr5dD6E3hQNLXBvZXYAxo4XrSIX6ysKSvZ/UUc6Eu
iIXclACSFhHUGIiEN4BuaFP7PH4PNc2Wfvc/krMnhFC4L96DRNwxF+4YrFclrmvdnCd4L3XpURFA
+DcXNUW7gOP8FOfEwuIS7c4eRFtNuRhYmzM3Zipan1wrHMww+LhNT187uFWTWm09z0vBMcubU9yB
iHoBcpEscCLUAElddI4XdD7ENDIgXJDu0+ZknkaVyoM2gD3tE23HQVT24u4XASmQndE+Mi0da+N7
gnu8vMYbxTrkhzeIrols8UezRe6dlQEJc9arj7MRydhPvWQNEY+lXdO+AjA8Xcn3oTxl5JZ4dJ2f
AL9B9MCK3f8hiYSXCaP5ukldCdkDt8swgQhkPzffklVoDyL1Dr157vMf3YIXA74bWcgFsWpqSyqX
Y1UvgzUXQJO4B30W3OcB9n46hL/ds5LxUuQV4+c/3r1dlVyK5+GrTmhPEjtnfPNd7txIbTXNtu8P
fayeVAgzlY02mCgVKM0xqdLSeb0OyN2SRBtCbVVewA761aJOaamF4d//KUN0OOdfyW6Nzs59GCPM
kaC0qWzUT6UVX6u9kQvLdALF0z7Sfar+crw1jaGfB4WEniTuqRK9+OFrzIvD0FlmobX+UOaBgvo3
0ayk15ztRGNIYjcsPrkk0UChJdZow4BHTgSIuVEUgjuQvAZjsfUTEh9gyp48yflhLkx/YD+9nDIo
Eyq3M2SDec2QP0n+H/GSW9icvFAU4gc/zB349O1QydK453blq/euQoJn5EzMPP21xQhGvuLOedNC
jtbrf2pMkGKMUgXWPTrOmbFA3MiKbKm2nU2uIN1n2+J1Ebe1pnb8abjD17SG4P1BNLB/mENuk4LA
TnQ6SmkBpziXGOfaPHQTXRroEySqPTGsuCoo9/uThgrpOGltXPOdG0T97NX65P1t+TOG30J1RLkl
d/4I1CQqAnB30xTs5l3K2gh2nbSbhz3cEJxPwti3bRGD5Or9/ZoyrEByyxQvxa/ISWr+qFsIqU4A
H6PPk07AcOL5xFPZpX6gH7vbv55fw+WXME2PESmGCej9vf+h5fBj9blmnA33uKE2CwA7SlUKqwhR
BHaBW7URt4LGX+vL8Vu+mFivD/U89sT/N54P2iNQ9iXbh2nxeiSSWUL+l/B18kJldJjCcWax/JI3
OivptHdbKORvoZWNNPRZIAmWVJMJgpjUIDUxY3RUA+brqjn5nx6kefsZCXwh+iv1Q1UKqjWWEWxO
QhDxhzz+YsKnEhbwolPhXaoPNM7UDJ8nXwcE8r9/NYkBjw6/mgK6m34UM4U/xM0lGWHmkumV8Exs
XeurRBbNmUdQpke1K6HQ2KkwdT+OlI/UxRF1Bq9kXlJslizjAPgtyc7xhvxbYjov81/Qbj98AhkB
7g2wtef0z65gcJJJxTswIFKqxmCd/e7Fr9LuudkGx5NiurpDekF3ZKsH+7viXIG4P2axEPd57k4Y
7iB54sS1NMfjt31duN3YWQOJF3/cpQ50UHc7IE6pYzLjV9Timsk5ppPIZ+qjniNMBP8j2XB7EQ1M
TqwQ/GWtiunO/KMKUR64Uv/5gFeU3VPXYnL2Totq1xc9QXy1M2pXWFr2qOhqEJwEXa8DdEpp25iV
9QRyKGyyaA3PwE3op00Rqxh1qhwuZ9mwpcZn6N+D6lI/mloOPfgu73HW7tEuCka7YS8R4a5JmX43
gk9y9q2j1CkIIarhcrMk1Pk3UsOS3gyQYCjh8nYO4ipl4/eRikr8Ip4cASbBghGDioxk4KzZqwI/
vM2uBU/dMRRZx7qvUI/F6+ulY2dQUOfUxdHiVLDWjkiVTsvaxFQoxoeU7c/2q706eFySuhRG2g0e
1bEdpdZEt3mUaODFDzZ8VteFBeYyn14DwiGHtzzuhVzFm1niQCwZYvxRDMKGfXgMB95DSQbFATae
pnL7gsGKkagAFrwq/OK93qUXNKD2YrW1V2rJMTlP/Rjl28shbhkhE4DU9fJs4tufy21l4yvvXp9r
W0H8o3BSlnRA018ljq6WuX3/tt7Kw+W5Nxl0smzQ4T8MAmtglt9cNZ+ZxpsRyb1xgNL349vJKdqD
CpU3vhCjBa3Li47SMCRLDBvc9ehejEy6UFcysytK7DNKyb6wTm1Tl2Hf0T19/Rm80bBBK8x4FH+2
fLF6yApBj63fGWl9lic5MX9Q2YFFt4hIMWYfOM2V+cyrAJB9b8h6a+LyvRr2DM7CDIxJCGg5zb6h
t1x04YUsBBROTUdZ6I+fQVKEQ7sAX8jXRxxkOm660VobIbntqiJ04T0+rCw5RRsMu5+1a44r730O
iSFHbO/runKdkIgBYIZXZyQr8vMXyi7YjCy0PemWhhWdsgRMF3xT0za3gy3g1jLNAvXcFw1e3Xpx
XNKe54J80UNWeJLBj440kABFEVsdjEWAuvz4dHPeKceLphdwPkesPvYDjObDalmj8TS+D9Z+yn7H
z/38CkYB5zHHzhANjToZn4blyR9zN/eYu5I5xu6QsJ+W1hVnz5j+I2NHTX7j/OE0Bu4chxnD6mtd
J0ao0WcC2kfBWQXoOu03tdboI+Ye2beLacnSIyLD9B81SH9YpBScDjkN+GvVaQOsWWeRwzPnOSiO
NqfrhWePkUqI6t7WT9b+9pYjfGN4/RR5gzL9yvi8oDV0hpv0eteGxDqcGN4YbEabti+cE6ZJxEhO
chl+s6WFh21y88qob/n5bagZLZfePV5cGPNIU1zBuNGAd7Z4s9FNpB4r8aUeqZ5M5XkXvmK4PYCC
Avqh74Rq0e2RW0RD3Qygyy4gio54TT8wBEB16rBjlODJdz/J9J1fpJoFAIg3FLjwKK64tnCEFQir
UmTur0gtD3osAaYoLhcJEfi03nV3q0mJTIaChaUGuH7uixJJxovNRXfIu20AeWu9IUjcSMlkasdy
z+BeKCImbVVzgBN8pbWnld5AP8yzEfs6wGas6D2B/R8aT27Dv1Y/ClFTcoWrCBMg4TAUB4k6ml2I
c6u7mn6Co1Sd+ZDBEgO0aMsy5lNV8ACiJs/SiQngHv8JcKxV1Igxa4luJD9hDGQU2buMmuI62e4M
uk0ijCUX+bpxl8bhgZ6aLrGa6rAt/hItWsXl4GYqCw07EK+73lO9PnSXlnhoDg2boapy9WaB2OWC
jPN4/9Y7ARI0PLoHMQNvfHwW3DbuMHXmeqMMo3Exy9ZEpvOQTnEB2/1zXnRhjEDYJzb6SLsBN6YG
q96G2+lGGpcq//o1bSmb0WABLdtDSxRqHf2r3O9scRTYNaegg8qK1PebT8wc4wbRis+LZWwAdsU0
XERe1nRRr+zqPyVeOnefc51xwOwBz97JS7rSrSnNF8pSMfsdcthHjzIRKv0ci/OXEwgsEZ/n+Z9W
SXTr79nH49bj2TsycB39MIYaG93ndnbLy//OvjXetYCOby49LmtaFtmXqNm8UX5pzKUCLBkihrZ1
Fuc6cVctmopw8Ec0yk9Kw5xTucFGM28rJwxqE0Sr7y7rlD3MH/21WDahU0hPH1GLgc3zOpDAHDsm
B4SjJ3WsTUx4RVveLloBG1hUbB4Mzoy75GPH8/aH3dD/nJXL1blFOE5j0xN8Bft7SP6IwRwbROOt
evaDu6Islhb4amSipwwI9QRyQUqKHVIUp3sslSMySErf3ggSgvzFL2tpsXXAKphm8CdxX79euNdT
feNjLG5xOLDBohFfzH8VecDs71gCeIktPhLdVvdTIoaYvU581vfiSiRG955qiJcnTamcF6hsREI+
lMFfU9me43f2SsXfuhXUB+WUgBXgGc2/Vvv7tNZH8noHKc2+PCxQ4m3gQDxofHgUKLMN9MfhkEbd
gzww0qQRyp506kuQ0wAMgosxcTiwaoU+xUJXEeQoZkNWW7ijkOWJ5DLkQI7KFfAbOQkp64LOYSNF
3xJhi9jquZy6fI4sXLtEtMc+X/e4gK+cmSB142A2+FiHNCcZMbrMMmBEq5tjpge4qIZgfSAPUknZ
daH7hl7ooHXpnOb2MaverRd0kQmFuq18pDYYBo0UP7Mm5z2rIgGXQQIZ29SpgrG8sDmjYRwNUlaE
gFODKZ2sEeZke5E0gcTTo14ct3yL52XrbrTYw4TGmqkRq3HIuWM3OOWz7wSs4uMVFEhSEHfR0QeP
EzJjOxunSwmP0uRtZxEusP24i9UvlTLWNfHKlYSiPMgXGvv+/zSkMSSKcxm2szxToAJKp4IU5Gla
Lk2G92oSFn98PvN+J+38BIrfNh0iGaQsVFIudU5z3G3moK5SWzx5ZcOIPvAkHTfsXAPEEdWQh+Ii
dn5ILuFm6SOUIoRf4pavsK66Gu+H7dRkekIZ9oZgzFooFOZx9puDz39aYpajyCwZfqTmkcGn4fB8
ln1g0oJneMKFzKIFs3WHFEVcHKKrQL/LXvVtwjhFFUF9QM4LpdDizdiRjhSdS8R6fcMARw/QtbL3
JgY+4o6EnOJWbyppHJJnsxy5N3T3+e6Z7qHwyVjMyfu1wOFT0hzeVLWPnCfDeGCqROLww/S7yBEs
vYK/XDVDoxVfPk0pO1CQsB49buDms+6S8vM0UGjXK35tVvx4DJUTKjw3ZkLQ93Bie66+LpMfT9je
ZYqbhB5cNmxB9IwXa6BwOZcEYow38dCvD4wLS1V0WEba9QUubVBrnmUala+uKhLUsu4iIE6xVsd+
SDfeU2hZxCbbAVf4K5GEXe+H5/nisSFm+fh9HvzPzMDBfdS9TejAaWMPeKSA9JdqLNdJDX4fZe5F
SjbUDUW9I3PYJXmhy64vu1DHH2yWATWD0xAgGzPfOXld/am726pQtHs8ugNr6T4xdgAE5c/CNVOQ
7Arzhtuw4m+SIh7ACwShxIzBu7/yIMNa1nFz5cK+bQCEAl8euWg+sNlbaxu+qQ4T4bPWK7RwnyNF
7LzMmZG2PGELxHX4OfP6PbRPab33YBjysR7LywWgSgLASuERAQODGebNYkhNnURgpKYMo7Q/4PKA
QrfMOSfnpPNhnITccjL88fQ+yV9PcO2LflCja+xCLjZ7mV66lfIxFzq5aAqjcfEIasCS9zO2ZwyX
bdxR6ZD1mmOV0f+aOupeWqNg0aCS8wieV1TU6Tvt0akVIPWhz+FXmAWKr4QI6rh5/QjOnRvUMhSi
J30JN6w1qcyBOlQywEeC++FrB6jaREQqabJJu+L/rNNWFDGI0Di+7Cj5YC+9ndXJSjMVOl2S+btU
waJZdA/zJ9/5pPbcxJ8pXPdM6gnsWe1wdOanwMM2FijfA0f7zG6z0lpByFz4g3C/koLKDKxzp+l2
l9iBqSCVyjQZnPFmXcw5Z++aQU2LLqAcpeoa5GZE1E2kCVbwk/0F+IJ1upteiEQSRv7PImop0XR/
S2JUDvik/Q9cofAsJ4UNP417vS9mQc9/00/rluX0c9TcJpq1QNv2GaT3Ejcw+2McEV+pmTFZxGdm
Gkq0WEizkU6+rvGmMzIF4YKe6m8zb2mZx+tuxXqEh/yT7HpAxL8OOdW9MEMxMM/xmJIkSKVQbURu
ofRUGnjwNgAhjbpzWQ+sQ10Dk9UEp6pl/KDJGbICLVlYZO+JCVhpDxBlgDxFONyQ8kdWo+WuFTgH
DL36XsYKzX9o66EQhmPYFNss7st4+u0mwQlq9b4SMijoMppOipwi4dveldlMS5u0pIBdrqZJSTFC
tpa+33MZi30eGzXEoAfg/bKkjsQTc99GHleZxsYUcKXFup3unBvW6qTkZi1IIz9o3qr2PMpYg9tb
yd/F2Z2KzRSNttaFXy7uYmfXRbVAqDAdKhT0/ZqaowOdouplscslD9wuLaJGrO9G+9z9N8YZ+AUv
9UMJBgPBhoOY+xXHIdLDsgEE47oHZryWTEq8DbkNXR+s2yT3JXj7RXwvJJLtfFqAMNUvHHyHxgcv
aF/j2AWeZOLf3N2Afp+cJWdS/sOBw2RAt9/iegryrSlW54YFuVQF33ls4Rumd7Rhxz92ODblhw/H
FnL9AtiGlNq2GH5HunszwFhPMNjMzh8o0dzcW0Jpwy3HcJwzdlR9OpPCc7m0bXr3SU1lS7C2J64c
XZS0PCozYhwvzaa6VWMNvOBon70qwe8WZnvuZFCxEog/dJ1e4vRXYcty4Q9e73qmg9JqW77Yo02o
UJaK4eZeJTG9mUrVu+ZRfInoF1KDbnLyeIfAXn/SrKGe/i6LlQPrxhGGrfHEvVxiPICD+U/yrmsi
c2OqzJzKfo9bDsOy0hz+WEH+yVmQYvosexA385iqm7anNII13MX8uLNPEay6JDGCJL/RDcHFM45p
+zeEmlapnd4UpWs769arU10hwk5V8z1BNsLqqh7C0xtm1kcK+EjAHxIZglhQZyijzB5m157d0uY0
Rage8aVnqL2UzMbe5E2Zk0npFOJa3MtTHGRRFC1/EQJjwRG+V+sr4Yy0YCgJ9cE3/DU2qGGuhMVx
HOmg8TwmHmK+SrWDxuTkzRfMw+CuDcVBbQd5Y9DZLyN7xXQEsveZMhpwGOx0C0W+uCElRVobnnIS
IgHaWnJDce8DxIs0jQolO+tsYBXWagIB+b1w2CfGRovzwDKclckBA3dZJehvEt8JEGa64nq99nSC
j5cuhyfHRkDkbWlhigqm/4BMkiaQFOuE25dGElLMaK4woH9M60KukGUxCsCKUtFmh/p03nWDnNf3
9aU/Ctd0OU90Sxea8vTGyESxOScFplSt1W3WwoyUUqFsodj5xrd4oxM8XnsPypoxrmu21SupIrM+
zUlYm5+dBakbsnt6iAUrDqwa9aUzkfL6OxjWDvoq+3+0eSfO1FSUaSpxTtrq/TeZjKCuc8jlkjQI
vxt6bohTcPO6DuQElSrtxRoAdI6JfIddusuR3qKQIr+8qrGl9t82sHsntP/u6B8EHtEQzbk4Dfks
BB0dFqNQCGUg0vBJAwygJ2goFSq1/lcbg4yM4tuh79lWrrFMn6PSjMrjhvIAytOCGNgfnW+yJ5Pu
c9XaOdcQTT3BYmgkAdhaHLJp0GLrxZo49ZgDSJbRJH8ZBnJKFiqJz6WWnaKSGM14oUVvlPWVKbXx
tpiabUZJ8Xead/fn74Th6RoCc0EweflnpslJ1ipFM4hwHDCjIQtKMCr9wMMbYKRPy9Xe60DxlyUq
eIo4YzD78iWmB1jpWMAA+2Q/eXuJOKeLmyUPn2z3rfKa5jXRw1auhs9qX3JVGAAeOeHdi74L2Lwr
FL0Suit/tOT+r8jTNnTFub/+qASZdmPXvxTezxl8JEju5cG7A+6Ch9uFA12JgxiZrh+I37Ft66mG
nFTvFC2pR5qkJ4VAO1KxNlwJhojIzHQbDb0F2RQMACGgYipOIMyaKGjPUXBVGTNbFUDpzgWsCORD
/fBbvzdhJB1ssqgeB6KuXbmMGDKkBqEQ2Ug+cVTV/JKkDHI6/zru0qHQoLgAc4oPbC715Gmc8V/9
+771X1KPuqb6yDVto70I1f7b6CvCWJRmeU3h2Q6PNegpOz8qF0o5+DGkuHtFZItBa04Dbb1hB7Ra
j4qKP7Eg6dwM6b96z/xwF/RwJMAR+7CYFiIaE6HCEwpLcQUEmQ84fQeuo3WZ/fk1FJDpMwrBcFOS
uyTLpRKR7NitnNSoN9amdPuxfkMWbLAtg9Z7Sq9+0VETRen0qxvDw09107s/QKzQPWYwoFW0NzWF
lb9tLUDCSUIzksYdm/tTYS334yL/9evpXg8qqQQp9GlP1Fe74GLrohCqoCSXlncRMKkQJhnn8b04
72nhFxPgisD2JlFU7pJWnVkLT65WhHsp5uD6CRrMNkMSKhAnmHqXedyuisArA5eIRu+UWwwx496Y
IukF68sUH3Ogaw3cCsx/ka/dmg3eZMxtdGSDuzgzg8EEUBFSz0Q9iNTQcm24Te97HH7i4GMilO/L
xixiiNL3kngl1m5Tr2bBd9dunxw/Y40gfZtgV0oUWiEu/Af6tqTJEhXr9ogU7ac3GMTsCZjmITvK
7ZLDx9sqdFPyzTAANN4o619Nuo65Jye0eiZDkVz9O3/Lsr5VbbVby1rMwzvIJbZixy5J4GAVCRXf
QuzpI3WFMxPEhblIBd3t7NRJQpxK/WnOqCusqGAXJeugUuy2m4SBDnr2/2OznNsd56UsX8PaW0Dg
2nkPUCLvsihASga8xcg5dIelC3NYRF/rfc0KC5q6q88Wjwb4E5GQDrfm3jgVJbGlQlfxQDUAOvEi
FFhVQBqFbZd6dz99SNh+OlH3gNAT1wm4IJHHrEZECBr5BygXAMZh7wlh6kXOUtVRgfT6f5ZGkNGP
mdRv3l+OXd+CmLW9SzHokbVJwS5D0cQpsFVRv2aYzl+EGASlC2sOD5jlEVuvvvtQIJrnZiZTpYif
PG8UoCSL3A1Bf0zYuvqNGoRayW+10m6MYVdfbWT+j4MRrH4ABdRo7z1ZAnMaT4+TNjg5px32Ajp8
xao3hI3QjJwjk895wRgZzLL2d3TloRkrxeVIUpDhryS/9w7011QwTPeRFXVEWlms48+5y2GIqYKd
fTc4ZCTvTpwfeZxT5U4mRbiEJ7UWvIcQg6SKy/wr2Fo9elx7YAAPV8qp6ED+vURZ8bzIywkfpv2V
RrXh4PZvEMp8Wtgtqkj9f32seBREaN66WzkBGxn+xaa6XOcw5E/PmSiZpoXCCemAlNktwaK4pyWP
7oBpad50yOig/UydN+ltPx2lHxd3w2YAPncU6S8jF1J7z6O3PlM7CNMlhEI7vVfSQDPLRKnQC3gY
mmchvbe7RO0GpJQWYvgYMZ0RJqKhKXJf0taUTMiTDUt1/+nkOxBAasAOyShjKAOw9qZrwbZjrdvC
lfEx8hxBvMmBn+wVFjAVS+9oos8s3YmEhZTzRMbQjcHYjl8JCC6gcf5ay1w1+jL4d6q5ry0G3VrT
mk1kchU7Hjj78PsQA3+g/KkTBJGW6QGIYWE58JCuFlO4eyBPnnFToJDbJjw9uNwRbWN4FY1wOVrB
HDocHJenvPzWevRxpcdJQlY7Uurosds747F091dIMVx15spMfMx8QfQOoEwHMSnIhCSTxuszDD3D
KFvVY/oS4qBW05hP+h2VoglloM3MfpswrzO2J/JiPfp3UWwwRRcrJHZ7JRB2yoCb9ZwGBk55BjD5
CU0n4IUyre+uz/fJl08/M0vyQfOSN8M0zJElsZlE+DzfM92DMZVD40ZsZnoPSwUb6bxAv0vX4+eD
sXCmCs3fQzr2XjVcbVEHTrJsIioM10WUxjYL43864+Z28+vpirRPt+ls93fzKUVbxIFrrbNHFpqU
DqPpjjBC4PRohdwEggWfRHsS6GVXgu6bLiOsylU6U4VxQpH0Bf4fRLi7odnXn+rgkhm8H/d4hh0O
K1YUAADyWqjyCqNoey6T02dXKU5lDq/rdV17jnQxTIaUeAUwO93qCxrWUwg/vaoSEtEN5fxqvoBc
CQykqfbRg+ghWSf1XQNjzcPgFe7bohxOrmjO9PGcErkowKteQDjd0KTQfMm0W/qLgsDVcx2BqKNb
qrrMYUg6iiL31F/lXEhuLbm3QWHJkEue9S0+8xB8bshcPFjID1soIo7Wp2YP2hN78T3l05OMbCco
3Yf7mijW6py+wdo81/HS1Fs1s11b1G90WWWul/c7Lc6m+wDSM+UkdmfVATIRLfRS58RxxME5jTq5
mQ7U7vrRZ7V4Ka84jcAgpphniGX+W873mQY/jUzNspRHbi0PTkyG15zW+5OJWU9GDF/INeLqrWMS
xW1tRei11fzddCNCVeyCY+LhTiMa5fqCcmt6QtdbS70D0m4XmCkUQbcSBM3xA+w313YiF3vdCMtL
ed8l7u5ZwbWLzS2zUpq1HWi/xgbtmsfm+dpIE6KOKJFYSvPNq1Q0gvZccZ4eMlDyJ+ZFkdl2rvN9
JsEQw3oguhNvtPlVH0ETyQlVN24vY61FjRZFzkfDGhc50ZN6sxBL01j3eSu4Pvjx76p6xBtNRWBb
zabjhpQdhYbdYp+9PwHiHxeHAptkDxJ5gaO1d3NuC1GWHNpM9nGQTB0N/6YzL9hDZEc2hgwF60fx
cc9Efte5D/96MMIF1zZXEscHwFENpy/IiF4hjSNsTg7WAWX0uT6WGdNilAJmjdVIG8zBouAXc4Sn
D6tkBBCXgbKvjcjmDvP5LBxzbqRzR4FdR5PA8Dt4U/8gYkU09RGuGALUR8q+jlQIYwor4E/pGhl7
RERR5Z7FBDSOVqAdze9tDsF+YAzxJ7hZqIa3/XzJwgSKHiwljHvNEgpxUAoMmkNZ0WjxnkiFc6Ff
31FfbWV0gK1tPADevQVYnOCH4SACDTcp6eHWMLNhU1mM1nffCG9D3K3YuxQDBXudVD2NE4Rn+VR5
mFaN/lGJ0Afe7gTLJdmWsQiPr2eIHevCAREsfx22nYy6ClqfGGpZfG5TmZtnYcukB0yd7VhM+66x
db7IfhWIVyamC92rmCrQeguEghwgdNUrplomrURlzXHwVLCSa7GUCP20T7QZwZnHAv6RZDZJx25B
BBqgrK5ZyKLwU5wkswM7x7Yzibf9M8Jw9ATYoCw26wLy7vKgOqR+CcAxAhmEAfbhvua9OxcUwdHd
JRwCzlJ28W4VxgYc+R7W+clcQzAAt/ePIk+Q+z1Cush1pcPb/ihhv7eBF9Nvyrgijxn+hb1q7uEP
zEVHFF1g4jQk49vRm8ipZ7nhVmf7+Bjzq/d8CkruWUk/YpXJVdUCLM1rSa3+MnI6s0xHCF8+vSDv
OoQz9Oyk9S0nbPTgDJ5xf9ur/yxqjJKVzMCA24XveSYG+5hETE8yplbLzIctDTB+MPmZj9BjiRL9
b6C5ZYYLFpYcZWxoc+iDT1YCNKIJMwXxWvnlfrqhzrpsfHdaCPcI24vcmLVqbp6njytZPogXxtVq
UkleYkAC2Ky8RLlFBx0gJS09K8o/Wsopq1VodjXceHuiPWBgwZu50lCkJ2TZOMc1Rlh1quCAX9s7
AIROJ9Cex6Pg2lF9tW75fU8l5w19xc6HHs3qZYnhTuR7EyEcrtLCSEZSnyYhi072fssT0jontiEy
85l7ctjKiv8iImi3gbVyINN5M5R6vHUsyNQE07H4p9EH09YWLqaT1KnmfsOxNQWt3fZPyc8iK/x0
xbeVzOpSwO3T7hd0NFzGBkZFppUG4b59haBkJgTLftJLKcBMrH2D7tzhEmLVxPCDi07jSysRfiuI
lmKCtNwZ04TTEYJ4EwrQmDdXl6aY82AiImDEavj93zsN8dkFTgVoN5mA43/78d5HV8Dx8MTCRtQ0
OSIhJYDOtuygEx/3AoDnWzYRc6ni2DSHsei+1SCgqQUn/7y3m52LQv+ck0vF+I+Bx2uoOECNRx7w
Vf+p+WS7McOwVeLo4jS5OHlMqNg6HNrXVPfiQ5XuKYI+59AFq/pm0kbl5AZ2byBoanxQ0RE6V6BH
f5Rb/10Tm/W0Ir9wqSkXZxE4kC8Gr+4hSLaPRxScPb90NTifBZd+DDnlAwqM/9M1PEt7O8+RxXqu
LbJ65mJykqfUM/KB0IvDs4NMtkE5AGZvSgEEjccQ5EhDDTMfg8wtcFjYqwFSdKj5P3L53tjKJFvu
qrgTJiFGKb++QTZ8jfonrdsU/xfPxwiYbst5650yfIZQsMcTI+L4eo6V8iO7JgleYYgtqXm/HY+T
RChPN1RH3n+Nzub9xG2fj6J9mdteHoaMS6bGKkoD42wCHkJewte0F+E47T/NS5j/2vtFhnZgsqKI
uigJzYhfBOJTOtrsjljXe7JOZ+Rpe1/TTR1mOwtDpP1KbNAr4CC/2JvM5yJ0SgLAu4M1MUznLKh1
/c6a1nVFC7nAfzYLWtuVJlUakR3iWndjvpaQOGeHC+HR+4v/Ed/jYFR7zPmdE92PtrjpDamOipEV
Uxw5uOGbRUQa0KrZjAgGWT+8J3dGeYlKuozh5DCnpirno63/lKXUgs4atHFV2bQLUZF3JsVCr0PW
JnfE2y7TDWSpcldPmEA4Lp2e8RZNWnRHCeU3d1rWmq3pOsBDcnrh9DCSLW9Trw5TkJEp1CLj5C4a
37ChJUxDo0qM6MzoK6WsxF88atVlq+WyYh1tVQwQqlyE/Z5dH+HoqnRz5uLXhNqx+w/DGkrl5YdX
IsnnGyqLvX2+zokp2AJe+Z0UKzntm64uIufxqcPvHi08B9mH7q7iHS6x0ZW0IinsW1442K92AOJa
NEgiUKO78EBsZsU7OX8c8BrSzO7godSrLYaBfIHUwYYwxqvZAcvmF19C2PLkXOEuLK9TBuFQURIJ
1TjvF3/Z/LAnfOELs5y6jLc52w0V7c0GUG53O3KC98RKUSeFbnAufNDhl4UbPasLuEgixdB8gUzE
yPyBF8j/OrUq1EmavpUh3Y3D/qL7+78Lg0JA/eydgJathLUWtlFc6uwAx3iKgiXqGLNib8jidbFR
bLgFalTbkUtTK9Uua2cT9WYSc4rrXhnoNgOa3U706BxgRSiKPweL1IlT24M6QlN1W3pMnLkLCxqj
EZKvFOEmBUDmt/q2bLHlwd7HvBB1HM9EpmI2q8T9erJJIY00+7sNAi4jNfGoUJEuJ7N8NQ3AtZ94
0KCNlpVM+82JLLihADh1PcGKiBBDNb7wzpo43ZdnnMXkdGB21S12HyCC8mG2Zn4JOG8de81Z8Mpk
ZgochFrdeOXtPPdxEVYYT2pW8bDz1BZ8gB5WwQcN9vSWtDE/+RWU6PrLDO5KycyivSioA7aPT10J
WnGnihNlbgd3U+wDmB3xf2BQRnhrngQvaVqrvig6sOag8ylcFdaQRVFAxeV/+0KgD5MhEWYeOo8t
Foya+aU++1jeBcFX1fdKPCPvNURApczG5T3ZLk+DOiQ/Y4/+vja+6A3XIdTBCZtZIolQQX4wdODf
CCCBGXp4IcRcl7CBJAeOAThycyupz3uDnEak9aQyou0xBkysAwgyuMLEcBDZ67QCFAJVXG3kkyA5
oW0bjtvp4jmZPzCCt8nJ2ZfjUda9kLtYXZ+feUq6kTQzuYheEir4e/qoyUJ4Qgi58fnFPUsNEbOq
j4XaayTsZMZauicXMxYOE5eN3UzPzjVnGJoHaN0GVvEN6huMrPVRQhjy32pbxw6mf1fnaEWSdMoE
KzNX8dPAXGyjSTszWDOloKusd66Qmwpkd9OpJCMewPYwm76KyXrwLO1zWDby7zjQpAzDLYKCUviE
xe+xwGIuCwXAy613+l+ybv4QFHZpQ7Vs2usoBX4Ry6HDAScabtDpo58t7piSSdt4aPta59D+LEnC
F5Kxv0ZDo15T/g6vqmOJqPYCEVeBPRtzjXZ/dNrJHL0OLSGy5qf+HJmkCbVGqPBQ9kLfu1SCL1M2
ED8rkfac+IPAoMqqp+fEVrM2yQWJuJX7F33ZXlUOBVMZ7LZ/3cQ/QHB+b8M0SROl/vroVA+Tw306
uDodyVEAM0F2Yx95j+syypROU3NH76smiSbti4nKbCt5I0gR7safw0mb80qUtSKR4YeB4HkGXtIH
odCR9/fthqiRt3i7UyC97fcTld51Vs5ChZmtG6o14dfDnVLlHzaiw+ps6WBEUuDs9w0g6v9okQ8j
krABenchCkTipYV+25LSznToVwi2P6rl5s2Kzaad9Jvp1XvQUzUdWWGeFJdlnEIS/fKfd300SmcH
J26kqD3g8wop9bf3TdFIbAStHhcTtifOCcIN1eEsQhesQ2wJIzQLOq4hzYt7UTnatQ54UR4MlNe+
0VhOUZ6HnLu+OgidoEmhERlw71Afd6a2fdkjQejfi4mbUOpGSRK71+NHlioabYYk4192x8Wum4t3
5G7C1nZNbpVxkn4MZFLg9WGbn7Bh4nybKKzlrKUKDyJgN9DuP+OgnEPsXoSsfvWMQ4oh/zPtj7fS
/BZti7HJ9meki6CpTOUDuCxXLoRfpOI/Bv9XMoDikkFNZ311IEZbVTYGyI8D8hYzwmksS6J1feS/
qO1Ibjf6O52ajMb7CHZBXhno5biv0gkXd3iZUXhxLvF5hCC0Arh9t3VrGo76GhL72plonUJH+o4c
bG/SklJFrNr0pY32LJAO7XcXDSCE5dd5e/o2hF2FsBKacYsvxYiSsgX2WTkn+BnMp+yhjEXDgGGH
ogMGr6r0tHVTuWkG1Hb2OfuRMF+GLebRtEX54/YF/GwF82uChrgrqWsCGj0AXWR/4/SNdrDIRFTa
LgY/6l8rFt79kD66iUXLMEThOgvcJ6W7E/FAzl5MT29MDe/5eN4NJd3rXaxFKU6a0fqvv6vV4rd8
k2vxC34MSwm6Lot6lZrPhbqJswFZ0wjbz+qhL9sfyyfG0tj+RsehiWh1tBJgH0qamw/2UF6+hhE+
sLrfmdku9YUEWmtbuPRYjkztoBIooNaVAsfBANxji6n/zBCoWcog7Lb6Bx//GXy8PU3INMZ2IVN0
ljSJ2AvyLEexWIlLhg/5Gk6o5/qwQBeMzrs7J50+jXl+W78IAnoGIUwt34vz2jdl/rzJsR+IMx4j
xLD5QQ6Z05fw1pm9k6Vt3f0GiEbSjrAlZLQ3RBDugMntJjGNa2hqPQRi7cOsY+ASwj2qLha6Ll9o
7sJqh3awVE8yfStb2egHoAmBfZ+le7cbQnsXPCqm5ZoZv6QFDElV0Q5v+913poNXjDhZ06Fip5Wr
XCi0Wl+wW3OmtBtzxOd/BBSDUHsCUTe2cjoqVb6P1pPnelMtXli3qT/vH3lLCH57mu52m3YbQ5oC
zuqkBYPosHbKeIYAf+cRhi0oHaPqdXeBkrZ4WcgMan3jgmORBCt3Q5j1nrc0K+fErplzDzKvFNst
XvUDERAmda7IaFosiqmJKhsogJ126zmOLni1dMBRZCsasX101S/ldX2bQ8g4wICM9Rmw5hV6YjQ9
rXy8dhPIzh9wsQr4xhd5exFDz4WBExLSqr+BGMgTaBlE2F5/hJcWVdAnrBGbxFH87CSB0PFSL8Zw
vkzPoirBKAp2MZlGhbqDFE+Vup81iG93ic36eGDnR+pGgyFD3lL8jWBvt4Pn1zLeKNmZbhrLVRKv
+LpDJehJT+obAbQdGoU2hf8DajTXTEI/Y+rihtd86wNpk5rfEL18hJ5PG9YP7qdwOozrc8tDB7Zl
sYf+SukGO7m6vEBZNPigrP+fkkGC7kRNEv8oUG1YKU7wiP33irMJUyflk07cGyGUooMkeKiy6beP
9Bu+AHyBPXkTElsS3lydza+kSqSpguzhqQMjwjm7SXTqNCoLBpc/3XyVcD0t2tltYVcXAccsegkK
OsNNLx0oi4TEQQZA9WeHuZJW688NJLIdLlyEgBMHr44tO+c5RKKckr//c5TmAjq+l803+u+m4yFf
9CrKdDyXPHhW4BAFLg742y1PD4cydP8J2DZEDPOzuI8BMTGsv/iQZO7Zy9c9OXNXvROXgwnJqp/u
5zaWw+6HwYbGbgkfZlx58D4qQS6BU+7q2oE/0izYEKOMOePkLheSA9G0Vq2ax5MxgtF+mC4whmlA
FMTtOQIMPihEY+hdzSql/gEk4PwFb5bwyyG7Ajib+y+i6Hxq4fw/+KDf/mq5lsymIYqZgczU743I
oVSNqcNAVgXvka9LQGoRPXD5XZ0Okfm3UzrmHZPeQ0hds2LnVrfrf0AkYYpxWmSBxirmX+ib8Iqm
xXNbpFvM0sXJG/KmEU+JNzfcNCTuFJn+/+UAye5uv9YBc3hmGgcpG8IxGL6fUg/lbQ4jdeb4d9xs
rAlqndHQ0afeU2bMJd/eHC8t/ZHu7hihrOQcsYWu4f+8AZJ38z9ynHTL0qfCSlnENgcPKfhCWi+0
EQolySzyHCtv5dMIbGmTpOhDdOm9AOgWKGWyV18ZbEx28r2ejBABkozaypht/fxPwV7QAaUuoH5U
cJAP0gol7UrW6ffdzKXJ8dbqsTB58BataDUvrY4H7Zy3690PsTTkkO0Mp2lK/mFpjtGMNb0/qSyU
9ATvtQ+TaP9C2KG8R8sMIJ1anMhNXjdEglvB5xX4TOoCJvF0Rp+cpzBShrhaxazIStoDhaxu/Jyo
SpWEiTUZ0zED8sKNnhyvXr06MV6kdj44uIqvdBCek5b2rTZ4RGoKu3NUJXfxo87Kyk3QkaZCmiSa
jaQ7QDopzkPwTd6W8Dw6PTLArxQ7FzdqsCqmMDi1copRZt7FnN4hR69jvLqrDm93nq82qddSPZ1O
MhTH91CNfe7CwKRShlER0vK7hEZIRe+HLEAk9MCdRhZzUXvQIY/j007EKoHKYDz/1LSrj6Qjh75K
lhsKGzaWpObl9YKQ6Xz1lAS32PCLaAKnSkb1JCiOOfxoftec5/W60ydtuE6yXrxjB4YQr+Y2ORLh
xTf9WjxK4QudrpnOuIiIXJKlnS4AVQQPVTC8FeBYjlW1wrWG3eXhbRIYcg8MZfA4dva4LKGRG9ja
94B+9e3aiJLdbfGd0+fMKC0JfmZLof/3oAiCisX2oOVqzVqyIrl/ziEx+floNOGeKgGtkyresED/
6P+G+/Xp0GY062mOu7ZxPuOaFPhCnmf81B1g3Y3YH6lbP38gStxcDbftPr8Ts9k4HXyLW7VTY7c0
26/KyvJKfhfiKa14fMKxUquhP8X/pLJ40sMp0T9srqrpym5Q2EOVPwe+DBrhvT2335t6ohGYJ1vo
ijz6jG3SuirIUyTOdCFx1X6aaCaSAl+9HN2+oadMSncnDlAMRrMMXDUtAJIN9dw6WQjHY2rvpda2
fwqZNXfdjTHYr2xpXST/ZU5HTya30kSrpfg0jfWe2h/MvdsT/zjRAs9GmE1IBsayBMakiPBwdcQ5
NLlVU/IdlNA43TCisVnxbtHjrBxceIVZ0cyKjuWZMnUkhhsQ8u6Ldp4mUIvjOqPNosjtL0DeKj2K
k21JGwqapvCOOTuMQmd537EMSLsJmE0jFY+JuGoXQTYSixOVu8ALfBIkJ61oIu+SnNDqJmMZwD4N
eLNyeqdEAeJ4N3SMQobOBxV0fzmDUBR2ZKvO35TKdIfcBnMxtCHHmJDcBLkdURkeGXIDwrRDUZC/
SRWFbmV8DSZCbmdGfgm3Drnqa9XovA2cI7TDWSv0Al5EVQ9nPV7PPOnghyELSafT8beDTfJf9CFF
AgB35zgKionhuNt83YkgOTuLWpV3RUE1A+hoFpZUrgj0acNixl/ZdwkbxSDVCvYvjtW2f1Zqaypg
7aqXfvzq5zn+36JfIOM/lAsC0kRj4ge61uoEgBTU+dSWzKmOQxpsbHy+pqe/YHg9XitKSCIGrXp1
EQiHFZHtlmHla0tJYd2m8LpJkwiiU7KRrjlLWa4Uf5+hlj3kYapOQpiT1NzZCrHhcFy6CxHL4XUY
z0hGZvbVs3lCMc6TMi/Gr5Z0vevulYiGpoK5gGUUAhxs9dfhJ4mw56pq1Hao0D6CuOUyADTBOFXW
RWXqc8yZLJ8JlefuMBvrEtNAxD/NrM+wgGn/IXZ6gKq0z9O3DdNgd6WLwHt1fIukHVCDCNjJRe7e
hg7nKKyEqheosbzaVK8NKQZDWfVibq3JYEpK6157ebMCXhsfSoHuTV76HIoeEkD48uO/NhaASINf
tB3louuXQEQMTtajmjyzDbx++z3E2gwP4Zed2/8tFw9T2rQ/ct1/Q5kH38J7BmFIJ755uYA3Inpe
dW0M7PMkeC32CHs7j938yBnI1vyzdHJP9UqeeFpHsrS9E6KKXjb92KZMK1Nqi4KwiPmkJD6epS3L
3Lia7TLWVqvrvTcXJa8E6ZSRfuqfYPDDtol97pmfXxHkhes+hrNmuSCPEEk8qM681h0hFYO8CFE6
ti+xTrjua1gScOuxJZez89GYLcL3SoUti5XK8NAoovOFJb0SVY+oVPnL3Re4bIRE2ciszEhWSgbW
4Ln8XZnmmu3TpDRXFR0pcqpL+s2kf6sx8vh8vlVZ32K3z1lM5pQuslGeAxGBoT+4ceyzZVglwgyV
v9T1pbOOB7txmuADyhQtiWmBSN3I1eJ7NPJxbynQ2qlVkl8GeUf3kS/fcKV0daKo2jMlqSGrrbUO
QvygoBXCDXHgmRisvQkzoY6ihBldayr6aej7u9xYgIoIX/FKSqXH1cnHg6tGkhJyphTu2C/goae/
ZCgamZHWA1gaLXY7OeZMy6z1G4MTNPVRMdKJotsawHXr5sMm+mwgjHRH8WRLbPcYkJDTOALd73VH
8iFtH9GC2mvpfVwUpdYwlyV6uwcCiqrFS/XhHbE82pxcEmqUHn5tzAlTnts0HNkBQDXab0LCJaRd
A7zPbht2RGFaZRO2SQ4JL/IDpGib9y5WJw127zNpu8b+Fwt7CNmfJn9q+Wjqlmh4v3odPAsRszIm
ndPa5s9PPLPqECjv00/RBDKvE3dlEhqB0/IPsY8vw2xF3cTYouxJq1h32W9RjIc1w1QGPe0a6CCa
YJR2bpg3+kWYjfxC20KtTvLrIXlH8FmvGbF+t7a35kki/7WDEUBA0qyQap1nC5aHBK6F2kXkaC0h
HJPeNqpxTgQyKFjfUCw6KraFQTPI7/dTjRs8hM19g10sTMJgKFOcQF++ou0xfZxpK8MHHftR+9Wq
LkuS25uxyW+BmjjCIozP/fPTzmD3A8H2D0+JfudoUAtx8YluRoigj6xVkj7mIvOyEF0XqCH9OG37
V6oSdfDBLvs3cBRFPoddWCgmpcZVCne3T1p3Up00u0HSm5eRrGO1C/IZ4nJvdo60nwXnkdSPojjX
eZlpr6KnNJGC04XtTg30owqeDOkgrwmsDpe6OTY94C6b+Xs3J4P6CYWViIh8JjfEpoUhJIDu9cye
oEWKPtydFyeeYbuZKcXJtr9/2IVTlVv6eMeJgDs+HyEiaBtpGwps4nAL8st6jjs/TGMNRaLrr8oS
w6+879YfHBk+tPR1YkPwGUUa00oJ1S2ue9GjXoI0CV3O1U+T8t2cWtV5TkPsZ9iI4v8hDiIqTEhQ
syCWTNRuqG+F8B1kN14Cdnp1sbTCZMsRQ2MUTUoV3G/khIFa+B1Qlwzdt6rKBQtEKRdkhw6yLiXc
Wy/FthwSdpqUaZd8bVRe5pASwcHXovQXOn78Nw3HX5Kz/DpKKqgrN7uR7kt4DynSDRTKfzOw7a4o
MArW1vM/d7dNSxvhbM6AzUVv8UVPwRwrtDZnWOeTYXBsbhs6+qtDMLxt/8e27umiv5xea0oC0rvd
okxsCnTgkVu6kRDfJENiSUVwr2EvQg5Fq1dhDlwobN/D6RvPktS4Ae9hRyNPdYFHglgsKf3sEPsa
l6QqTVLGx+o6T2K7oCCa40Mv+1TOnsS11QY7WImNE0um4G3vnDAIAO62aJ1s60If0F96KoqT8b04
d0B0UJi3nGO4hsRgvy59D2B2IwsiOJw/3uZe4Nk4vyAdBSVUSMmBHnJaJGYuBTOGSVzBX3G2whMd
ysSIIPEyyah7Gshz4WGh/E6XC11xI9vEI/QTW+aM0QxbeCLMXSaHZ2lJMUCrWYd1RZ7DzvnD4nGg
jyH6h8yQvpiwJC3kBpLndL3OmoI/hwMdtS/VVmRMfvaTAdBQ5eLmQg8fyvLrLAJlxDrn1QXYBjhf
CwpGWzdG2KQeEUY1IPc1L7huufyLaAoJmN/WxqsjzCW5Yt0MdL9naM1Rd9+ieZpfLiLQOlTPFMQG
8RY2CR5DRfuTE6GhT1yDFfHzqj+xtbve7MQ2apfbSHpTaGxbpAgIeJqBXQ+u5wfrK9Hjj2z4iLT4
0yL24YZm7x4LaURlvLkkRpEHiMjFcfsy6R84S791Ucy3WhM6KiIPSKM0XXQybXbhNWzNQMB5QqB+
RR0H69BEqIsKnIT6Kgr70FSGJVNTAhfeGk6RAw22DfzjZVTtABKKNiY3A0q9Br6z77GIncBmNMw1
FiKZRU9H4DXmJtwL3ZRiGEfZ7XtJ3ZU7vrckC5bj81HPWvNfseg7u1s0zY6oH5Yp8tq3cLx12SJ6
615xKXi0eFytgPu8blm35O8OD1yKstvoOlrE+Ylue7IwXRqz5iS+66vdSNfjUwiADpuCg7Jqm1Eb
19TIh3JKT/baj1qm/V72UqPpaUqsXG9epMH3Ccm50jxoCH4jBzE+5Ra9hw9DazCBzkJaALzIBkU/
oTfp4XbS3nEbExQE5JcOcNeNC1PTxOqtVQWkZSne//3+tK0dwIZXYtOfoaM1RCaYCIRgAclczxAM
nwu6S+OEJ7NxYBuc6ANIZc2c1FH8igJ0O00BMsER9+7IOKhSUTPjyLsZ1/Ze7qjDaNYQDwEonyyK
Ghv2mRifv9hS/vwy6JazpVL13SNsL5v4vRNGgexVbtNRkLe2PT2JtW/Ogdln6jYK5dpfQ13PHiVS
nifrkFpI9MpxiOQaEER1h8Is7oRgClxIFxWN+7o/vxwWEBNlBdzapoE/x4wGHiYKg55uM/7EQYao
OL813ersl3co3AN7VUp/6Us9jGKnjgiBiXpnlEgvPwVtFXbQyODP2dkdBAqxXdUrx9FuHsOJqPkN
3dukUoh2XPi+ed34RDTiekLxcWjxSNBJMLUeGw85fLIV1ygwoRTT/7I76EcQlZRhZ3iIbGbpHlYs
YamHilXloQ/vXe0ISs1yLlfU0to+8/tZCBH1XcJGb6PiaTvB/LDsjWm76RbP6vkQHxWUZcxnHEc4
RX2SqEYQOUycwsssKvOwMEq0qF+ESgdbWRHRNVjXBmu63I6mZsKwttB4KH3BO7Kbc15AavBefwkz
tb2SrZUFMR9MIi5jIVpQDGxuSwKXkefk1C8NneE8s576igyjjJ+zXLMpXhAOmqbtm9ZdHmAXRpdg
38WpNHf/l+r79k1tmJSGxHhuJA1dozSGsEuRsH/5iniW6Egq4DTeJDztq8INH0kbPmlN1pa4BEOo
IrBcaKZUpOTnJjq/DOsVicVCveVBmNyC8b2DzxKVLh8M8l6RU7jqXknECfTNFeXw6XyzVRIE+ULL
61whYsJvdFEQ23oq0r5IXd9O5ssgHthIj5ryEWvoF43fw1tu8mpX+vPdkCXeUrudEf9NmHv83Ads
BVX6v4BxIwZfFY5WWToqAuBvbWJN/e0xDv5/sY5sZ0oaNz44BwG49zkiTPATtazSOQ/ixEX8odxS
DPRvO2USk7P0KlUPpa+OQ18kp2orIl4Pxj/9VdoXtod4yTPUs+BcHOBNs8y2nheqORuu3viXf6Z5
LvmLfom7lHxE60NiXLTnRTf4KNdaPVut7Yyzmzfqc6yPOfaA8fmFF/y/bv/9inYR3dEpTM4ddAhq
cEcB174ZNLinTMSO2wFhuxpvl6NrorALWuX6JFZMuK4CC7gaDnQByyxq4NUOBMRCfVt/0WhMJIeq
maeGraVo7OiKu8QFbNvfNP3ObkW1yIorD/s4gpmU6JXp1EVmhhaxhYPUMyqiaWzDcbGDvqiWVGai
a2yeqgTWXOrfzkssEIdheQWL3SZFgBt2I/0/W/ffu5wS9LfVOpgKy3C1foL2jU1qLVgfM4uRNXNh
IPonl0V91IApDtDWs2XzVqB1gRxSi4nfH15YH0/KzEewBk8/yjTdn4fGVp7W74ae4Loo3VoZCmto
/IRuVg4n742n97M4n/pl9jNYNd7x3LMMYlLD0qQ+bBGy3wX3MpxEjThFLb6nUQp0O43wS41S2aji
yq3LbYgDArw3w+Iho4WvH4/rLFAsesJuDnxpIG72oybU0rRFmNWPEBf13ZXmkz8mJd7bN9oMuaRp
nVuiGIDHAhRhVs7t3ybJmAO2sAPLL4x5EJQHpZhp6CHavtqOP2wEHuPqanRH6TpGBZ7NgT2/GOMn
OPfcI7OX18qNMI5weC+3N/hf5HcBQoehKwubrSfgqQZ3WAXEjJ+QUWo8FhFXMIZ0GtNDkdmJFoHX
HiSXab5t1eqECVUTpoX7geIJMb+Ujyj+lMWe8wAHs9aq0HrK46PfDRQIuv2gLwcChdmbmFDbh53A
PzEgCqU2NH0RgGpgRqXX+QR7QBmSgV6GsZwayMjprsFhBmwNXxPsofJ54rqMxraSlBi6939Jnbdj
8oq8pRrNfaz9do3vkLGnPvN2U4JNpVE1Li4n9aGHG4ExcAapKqMOijRyGPe7sZjIbl/1ESGKue4y
r5uY2Zt6F7N3A0XX/ajRJg4XNYm9YwdmUCrF6zASpIHi/QFZpQRcEbgCtDn3q/eVetFPgZw2l7Pd
h1ouji8oBA5nCvoen3gcgKZJu2YOOCArXial9TZk2A451ZkrZX1ONoukuE4Gz9OZd6G9XH2vn2o7
IwHKCDhJHq/Yi/Usf+sRi09qXiadFB4xc9mCv2fjMWUh5pfRYAY/vh8vPIsh7QdSBdCaECy8//Pi
/1rE+CW7SSYfJOyUMnv0N1xZJ8IlLn1217Y3ZewWlHUfVRFOZ50KB+pP3bg07WK+pp8RbW53IOLc
rSdrFHBV/IX+rUOwObf6HF2+5zlF1GLZuw3Xs/FQxVqpD0dEyHGc6Qx8gFpYeyLAF5fzibd0VYYu
z/pVqorxo4COgiq2oOxaXtjlLxmCbMhJzbXgKfDal55pmdaPKMdLeDoV+MFSrHZwooPuStr1flFj
6ava759FhycinFXvlFvD44HaWiaZBJAWeLy9vJseop1yCZAAu1VTCJ3rY6WK0eZ3pUpYqXSV9qdL
5Mf9R8sKGX3TquU0siGtLzJyrQkzMhFzhXSVN7p39cYoe6gj3jTNHECCuFMYlM6DFrX0H40cCK/A
YVADKniUVQL5rlQkOskCKA1bsUDbEzBPecl254UFTlaEabdcAsLJ9GImeauywwxaH1yCg4O6mxty
hyAhUXI46x6VLTPUfvAuQbJeB6qafr71CjVh9+XkSBDY/TfrBhhdm90IMkEg79/Mu/jetqZ19/Ru
Z+r34ChGx+0bK0MONlWIN6SVf8yFrQVCCzGH3XYDM1fSVhKUa5oyy2D2qk7yEIwOgoUYV6OUBVFw
Ka+VeQ7stZWN4ucRf65hnuVyaK0e/Jiwu9fQ5Cyh8c8HiwpBYVTq7Num16jOE/GT3LY7MG0zZko+
RdzPvWc4qIWJUSzDlHMUpTi21H52/5p4uwKQUA3crjHiEsZUW/6Iwp+yKhJX09jpIWmLJXWMDdGM
49SnHdA2YF9FPIqGnK8UGNOWhrerxrNUrwM4GLFz+VuG2ovnzRuTXYOxxj90qEAyUm10olz0FKFg
z/c/cglybucQuJ1vhf30tvpbPi4jgtAeVPOeuyqUq5WR+SA7s1noOwTTWjpzGsoeyqvzvTZNx79G
jClPdAu/4oNlVh/Wtn3JUNp2D3XTDqFFjBgMa/pmJYqQRD0mHGs6HreA/n4/7kKMTJ03f1/B3WlW
jreLQaWO6MqzB59kf4hqNgUdF6l358Qc2g3VZS5o81J4se80eueOMQR/e1/QPVlkIp1pKeFJtWLh
MIcmz8+XX9lrCNj7LZB7+LqTU84KZsoT94co14HXlbNGV9HhBPDA+SNGYZuoN2JcRduo82vtKaHl
L+h2YoX85BypEBRRolD51g4AHL1u9wyntqNjwNbfLQRwcLQ933O6/LgyRbciubMnJ/AFSvRdPP6E
Q5aiN3nTVvlH+Z9/f2q893hBZTAX1BrsJ+iLv71YL012Zc7UY9SOYdkB2jRgpnZoxiO5QMabUv+4
XhkwLSWE+rFWwRCFkZWYQAvLOpVJkpAJvrhhH2nfmTq/aDJ8SLisqebeoP2J6SoS/ypqRwisKw0z
lpzVDYVff6PQ1sYCjqQLmXwpQOmneg4UEFmrDAH7MajTept+53p5nFmC3LNNxRWjTTKNGnx7kS0J
MjCLOsgCs3cHHbZK9K/Uj5CTjEHaEUgo3dkV/g7Y2Et7VOdXo8Un3+Uo1+xlrdKfO6q5YM+5f1GM
p8haI6gqGeL7+ArtNz/tvSg7M6gjy2IYq2TumhGppkKipzr7QzlDUlQshCeIBa6f0A4Sb8autwbb
6T8oGCKi+nuv1BAsIICETLDf9ICr2+IqPnFyQt6vK94Mp0fWWhjLgU14rVL1HcfgmclbSTH+Ri1C
Vad80/eG3OCu+H1pfXvk2twEQiZvm83Lc6GfDxhDnPocg3Vc2ofEBTuqWTid2i2f9vVhROSdlL06
U3d3SZWf0a6SxsauRi/a8etHGzrZJXZlfNXKbDalyHV6lxjoBLYTCubVu3ruqRS5ly3/kXnmtBeW
IxmNTjTrCY7ZP4WqLiRp/pspqlObitLPZlRrr+iuk8HwJinCUsya++MTiWral0wtgZ3Mxn10/hUt
FRBJ6OPZs4rXBGF3vtjw2YQK6CWDdDajr+p0/asHIR8GKvfFwwxy1p9/hZSffPSCDjax1LYPGMjR
i/UatwZFwiKR/NfyE5rBpyHyjCwIoLoJmMxoBlSCFFuDTsHatUbX175H8OENPEhEPrEFQLRA5Mwo
+oy9UyEJFECrcEBolXG3Jhhvpcj/Vrq/lBIPNNFqd3UpTTwR8WEpwBKm2O5dNRKj05amIAV5C3+2
OzaIyL0aM0oxUn0MMFQrIKxKqruFrhnZPUQfvHNUfymXP1Ig9TW/BMBaRWOTcN8Q7Dd9JwZ01lLH
JyXgP/vYjGC+qwF8QdGo+W6WfoBEsTCzdEjbxwmwy3voS7bdjIKlfKeuTR9iHkOwNV0nNa68IFnj
Y9qIcZPOSHT+o+k02GxSj4AET3o38LaTVeZhv/ntOhB4mJS8oBf4OIeLUbNiaBwYnjdod3mOQkUe
SBHahU8spOwM7ZfXLr+2/8iapmxpH1+9yC6FHmM4FzTk1mZcNTU955EjMdRs3eQBXZQ0DgY0d8NA
iJdN29x2kkiIFzXEGaPQRA8qdmyANqANQS5oPbCtL0A10siJ5jEhw2shnfZ+2eVSnp70zHOvRtDu
WjG0OeKzLlLRs9CsazQc6DMVimFpk4WGgXz3W51Jg1UhtkgySVoYmpDPnLwuN0AX81CfMmUL3ql8
yOdd+LXzj9UwG4IDksRyFFX9SH0sLIg9BWeJH9Z4O1ztnqyazy1RNXBqSwEMhkoADRQwzWc+oHfg
SOrQ6cKlZ7i80CwwaGJYHkTK14dVcI0/n+AD7eHS/4BUEa10QkEmSFle38lP8xJW3IX6rP1aqDIt
KPmflvr/SvPdLTKiCokCFWb7HBuk7QwNUil3nWcObyBigqtcGOweBaElBc+0Ck1xYgz8UZ1UAZHq
kxgrhrfKXEkzSYdGhIj4/6n+qkNmy78EtFxiOKFEyVk9WsSn31ToNpN5yZXrgM7xMEI/9zmPHz8K
c6wn2PBosF2cm1anehYmzZjienFLhDZ0jVCpkYH1V4JogjSb3Nsd1BsT7Yboe2DVjtoP3R7UgKOI
yPDg/T2uGnD2ZO/4r0cvRpRxqhcomF61kDhkk2f5pW7L2ta7kUkpTjEx5DgbS4qSjgLbNvTPRSpJ
cr37oBsAw2tl3FLB/4XspgenH3KILsRhcIWejFKUT1k755DsFuzaJnESBNl2+h/cI2J7BcN2oRgx
7hwmgVhBRU8m2KgiGcK8JIFt6ZzIKYLUGyo6v1580YBvkbF8P5TXuufgCrGDc9jtvq06xISRqvCk
87jx2I1t8I3NVlG0dhq1dGhC3UHyrmMatMrj2vnNbltu29P2e0xGi4twBaJ6yNjlPA17D8N/5oOT
Q5kiVBuZXcyf1XEoQQWQhwukIl2TWY/GoJ2alQTguOB7TCJXxjfmlTuDVK78AM37eMD8CvjKp4mk
wbQxIOz+4uRK6VE9YRuBdLxCld7iYX364Ce/AMFpSmHvfJXS35glAMPUyHr2QYElfPdJAJpGeXmY
KJOu/2wb9ABfakWSOLd5aYoi0/JlJkOF0lNufKqLS8vuI5lNc0ZVUrp/hLi8Qs7gLJ7SOWiBBd/N
L1idTRAAxN/sdcqKmVDQ8R+F56r+TYILx2QMJOsD4zJWizaakPLTMQEQNBJ0pGP8haD8J9DhFCJ/
Y2VS23ZxT0MmQOjwgfYzvnnIQLzkfnHDMr3nZPnhcHwsu+sTvsAW4/R2VrLod63Gzpb6xtCVINXJ
ayU5etBZqhw3j3t4fqRAJUP5ByuVpf1swUlbeSl/1UerHM+aPmuAA3Dy/qXFm3CemS3Uwig21Nmv
xtKZIurE5vMcaTGKDyReztYJdaHaokTuxwWbFvvXIbsN5CJ0/MagmrwsLTzW3COXw30WonsSZeh2
CEE0hoi9wKidlCp0YsxQLVNsA2MgBN0yzyVYCElvu0T0Xc7tW+/t4Pu/yIPdzeHv6nDnvhl29UZT
BcjCGZCqIBTUdqW14Ryf6cBZQ8/GF6ZNkD8s1ww7MPLFOValpfa0z9xkiob1HyLegjTGqgT25bka
2gVZZSLRahVgeOIeHMG0KEXZB9Pi5iVf6y+iyE0J/n9wk8Tw0iacXPHfDLlK6oQ9vX7VhR2YIgjj
wCkdJQhlY7akE73U9ArfLge7atv/7Nth6KWxcg1FPq2thBFh6+MdfKjnkYjrkuU/q5DkDLpSiiRh
BDXyqJZZXEhBx8otzv5ASxwLCUY+2htlknM8rcd8B8OaBDOECEef+z6NHKlcH7hXVzvndQvi6jO/
fXIEsUc4YJiUQShWyfFjcgC1MTaas0CLjEvMZC7b/J5ethBbrz4DNTiAtAbtomhHX1VirdtUO2oH
MUlArhlQcNGjE+giY1KbTL3uvorxfpZtaB/+9Uowa1mVtOzwYOPLpERWyi2ph06HswWVKfERcZML
Fk4Srj7Cq2ZjHX9IHeEX5O6WjlFuM1/juLeDqZwohNxjt7zCuXG8Z58vJsSspwQhedOA7rWQrOu0
QuRD6NmzMXQvTErkIcyRRo83Xn9FLTuCOoX4e9Dmno7QIteHhLG8gBSDvN7ixSGSM4vmqvZEe88z
lxOb7ysEsVFUnI6TZkcDG7vs3taL7AWuUGr3DDmZEAyUVmwCImPsqqita8PV69wVVgowTncLDC+A
jhdDKQ17eHCADc1xmoPeLEQwbhxaHo8laK0dzzbuHfez2pJtCx/e/dhL0fEhd6Q32+scOizJAQSz
GKT+hITvnlMR6gOMmwmg/uvI13TVMMATMu6T7fDRjwQt9//IrCLcLfzsVkj3E2x8qU/0lVDDB2bV
YrGoB/j+93Q/I67nWNnLX19XNjVTMl9iSl/SqSi8PPGgrjMHmgTeDpLEBVHtx90spF6x2A6xumCs
rMTapzOgcscX9yCQBq0b/eo23JkYiNA8tOev/a+2JPSqqaXvCuNsguafFNABIS9AWcTPtU5i1dps
8szVQI78CuEA4Form4IuZIgqlbjJRjmwMwi5N45nycLZ+rb4wAwLPo6JeyRrO/Q6bvcZQPEPWPQT
1MIjXHnA4qFFkMVAYuUNFbA6hHkcGGJ8Ixs0/HO+VVXCEvuo8cwB0ECutus4dwbEi7TWS3alx+vZ
Ya7L9NuXww4ZATCt8s0A/FNfMorEZYIeOjNR3mrM9/IBtETQw01jY7C1WshfcWDTpPxPh08lKnii
IA8O/yGg83v85rFOa0wFSNiOCpKZxDzA/uFITZ0fjSp+MphpL64lh7KxZs7K2M3yvjpdNCHbh9s2
77LwyEjhoI3gwA9Kd58iRBP8jknn0GoKVtC2DTZinWfydh6yDQwjLKjU7Px/dXPHRX7AKWkte/gz
/USCgMTH1Dyn6LI6dJeWMefgO4fxrwuVMIm1Ovm4dMbRz/Fl36RydFaUCVOM3I1L6TAmSkxw0G2z
GgA879ssB64iK6DMBeqLUA042NZINLsWh2kag1aFREno8nyPFIF31Z8KZFizA0t9Tf6ivcrawU63
7g1gJl+FT69SG4p6Dw+rWOVw/IKew9cc6zAJ2cUjW2DZidThXpXyT2bYKLnAKGmjgn2mkRUyVB+T
jXOVjGS8i/AJuVdUN0YTYqIXITNSeHMOpL+i/JGCdNpKIjxJ68FSZ98610vaKqPB0lCeBae9D3Ey
isb3soBj1UVi1hkhTGIBXqFNICQeJLk4d9iuE39MXVIuT2YFqpKQozG54MZ4XXZu3uJ6qZx3ez4C
ecUF9SQBVswKwLmCfCrLfFDQN0FNSZIKW0A6FtGFuydBve/EgvCpR4SaeCSPLe8zp8snSDsEH6hM
sZE2lfRd6AT+OY/SJZZ4UI4DOXeVfSTxib9tivPDrC3+QkDR6FwcqxzO2CSmJfABCSi3MM2ZIIwy
g0w/HypBoML6guE5W/VigNiPK8LnpaF6LYZEyVz4fj3D3NsOZJapcsIRjtAoCahx7KkT/N1TJY/t
z4iYpIVk5urz0dmI+T4Vg5AH3UpbJ6c6pIMDh4DW+A7d4tI+GjLi147/kB1wwbOT/2C21o+JD8b1
dZqln5eHSWADqyuGyFSh0czaeaABgxdhdr5aEdAzPdyHLaND9hkW36AgKQGENAXJq/0hBJ/aXky9
HPJ2UqqhqNGgQjMlYjdfKLlplVJhCxhhaWLfxVceLxEDrl/l265YVB9wyMQ7wbR3gkSSjhrLh069
l/Oojma06FPAN8ik3X2o+hqRqqL6wdO76Zx9/l6poAHEAE2SwgjnJBRt1OqnGpwNMGP6hh4iSd58
gGKracMvGT3MuKfWt2NLepecsyxbRd7U83ovug+cHdBAnGUPsWrzUeNHAnXdkQqm7KultrzuEodU
d9ApQK0cG0Mh6iXnKzY9wKcl6xkJflppBVbZFfl90IOGrdUAWea91Oe33TNFFabnWWpA7q+V/K5V
FX/0jP4f3JGNp9t6SPeru/0o0ngbp/dWr1Kalhw1iBH6nn+nD/mk/QrKwGebxyEscrEVvjOragNS
FqFoQQzQO+zBjBRniw3/jS7zQHR3jbxA/6JO1hGSUtGAHK6XTI+I9C1gRN4xfNwOzEA1kZ8+pnXG
jQiIM5coY3sSEY6mLa8lJOF+wAmueHWuG0ZdS6PSMpNjewR+d+oYxWJW4cxYOPEIfYyWCEJ8eaH9
JALm10jCga6ZuPpxfXWZykEzeAjpxw+e3QcC4HK/0NOtefx78S8aExZP+5YzofHW31ZrpKL3qGvj
USa+wQY6zuvTFOn4DTbNu2xJGT+5QrywbzKoUY0X03sSN10AilHgy/4e4qbdjciuo1l3RwfhMp5v
N/RdCp/DFfg0y57fJ1H0uPNbuEZRlKjLqbfeJGmTRqdXiC3lSZrZ5camhuXKClYvjfz/MuV3YNlZ
lpiC4++pL3djWRPPqLUULxZE9ATiL37RuC2ByMM765ISiBYl2lB+s+9kE/hXvzwMXO/vqfVYwn1p
21xveV8qSVVFf5Y3pGpeDIAACvhNtops97HDHilAdxbYU9x7KBxjMUfVdZSwMDTA7piml6SqMPtC
3JnE6NBCD33ryeP/opVmo22T+mAIYQ6GZ3GMjw0KMu1cooEr5o8cfZ8vzFAg+cZKyzGarkeeg3Xl
7ZagTT6f9HOEVIbd5P154ysmUXooKZLZjKxM3kY19zHykSB5kUWnwmX4k9cNWRwUGi4q3Au4R+hH
dmvNKpxL90Eo5yJP2T7jUkopokwe5oXliaCTRAXGwpTx7jiecoNlqlOP5K5LVkE7ypCFwMykKY44
3S4ds7E20HX+2BGw9DiAGwSELbKBJwvrFTeNg8anEVxsHeKBavqylLmWV/VYme6SmRBdUoMdqEkp
g3SdQRTPGYYIbvcpHE7sgx8CgfHsVPbKxeZvGUwjhIRUiCSBwGbM0guv8e5QBjw7AeugKPWW3wVz
e7HF3xE2sJewZwfh5u9Bptegu8ojOM8fQdyCW/0Xi0j3HxfKa8/0xUcN0SbPpM6FWeLWcJ4Aw/a5
3S6ULxaxkC6sMmwSwSnOuts4/OuLluczkCT3qttu9zGlkhDXDAAgNplYY6LWWcT7oiLFowUJ3DbG
eLdFOFyRqpq6OcJK60MeBuQwB4IaDzI20jONVJxTkUj9Q4nRzukAyB4bTFWS5UDzq2nueLhp3OB4
uGo+B6G6lVIFEgQExD6Z2FnaWEzbCQ2SlsTw8/AOxZeR2f/InWhC2Ha90dVUjYLeXj3HrB4QKxL4
/XFP2l3gUwfNnWY6I5C90PbkoGgw4uOqn+7lyBXq9vqCPAHBWXb8a0VTcLhDWOugm7c6aLhy9lkr
a3+s+HEAOpL9yERWhV7NkaqMbA9f7uKeAdv3F5NtCdCCfAXu5Am7uXYe8u3VLeJrml3Wb3dMhTz7
2BrLoJUIlI8L5W3W/rwpoXLlfpk8qPosatXK0LWtUzKzh+wBEYW6sA95oVUUNAt8Lr7gh66N1Kyv
C7ZU07Ks7k3qbaNgtpXWG5ItV10BRsldSUbJ2SVZd5XeDgOLuDBxPDuSL2fCmh8OjfW5zVQ2/oGW
pFnCRLJ8eALm5NoDZs8SxT7/xtRVqWy/2D8i1jOoyVpe5+dF0YcMovPA7Ik9hjB4hLOGCUMKm9Ji
1ZCOFqPRUNi2SjVtJG1pzreeoL9CLY0892UMT27FYWM9Y1r1DhWrGl+5lPjaPFoEKLfoCAoH2HK2
hpB+7ZpuEBtDukjBNL2YKoKIsiTfReDsa6kh9g4zov7WZdgQCjMCvgnKnK5wxYA7KSUFN9AJgp06
/GKE4X8QwDel8FO+093D/hwcsTIp2ssv+imbLIenKE3gOeC0gsU+1EBWkTHG1nwkN9oHtxW0bO31
uk4EnTtNNzwHLLCJEm2RMvwGI8DZsBHhcLLXYp2TRxekeppLGH9Eiog+OuqXyPyvhgBzlfPuAgBN
JVd6YMeiYQH7P/IgT6GPSzc6NsZyLH+htMgix5Dp3JTkdLG8SdCVwlHOdz/amtzdgPmBETfKX8Jl
EecKNXyImH3lc9Ss8owjMewDjAACMjOTXJIg0XqZu5/SBijqARnVgQWiVZQrJnC+KChDK42SEFE5
ZgMJdpkbwXrZFJNBmbsRBBESXe9xfyp58IzvtMEi4peM1/rDwzgsbBDxzZ1eScS2HfQdOjcedkf+
1qLIKwr4S11X0XDRvIvT7CWmimzR+g3OtqxnnADIYStoa3x4IBnWGej8gYrPSE5YM0Q4pAhzVS1A
RkmOKPJ+atW9Eels5cbn1BDlZgy0gAKRnAfwJKQyUKt8NPoPWD49PrZ+SvgpLIgJzFCNSboLQGZC
lwDLCzsnunOY4m55JyZMEgtalneeETbMZxQif/brNFTCbBuhzF5CBUxDVZO4iwEZyojpJPmyZ24W
sRndGIEJmhj2hzUzYedqY0nzBBivknpnZ0gTRAEluoAUQYUAeGZ8AVeFz/yyljXzoi3mP+hxafgP
kQ4EeFbMxDL+D3lv8WYNgQbrlsi64aHXxqnfZhf90VJleqxd5ThQAUs7LbYoeub9DEI5rAJyO+Mi
dujTntKyR0+pZiuhi6l64eS3+yU/KBd7GQO90FW6rktAlHiDD1Hi8n0NeaQQEpG1xyASF51xV+eT
AAWg6Bp9/LiBX8eZduQ/Tv9V70j0L+sMLkcCdM6onzhZrpysLRmq5yagg/4k1H2WM3Y8FLPZMuVS
ulFYLWKxuAks1RxUNUELcldsF++gdgSZFmO5TFvNqPE6xBVjiYTbco8Ix19+9eXqY3jd3rXWhbvN
+lAsyOfeze/3tKNYwqyb6mLjw+WjWiBJe96kd8JSrp5ZH57vLY1neW05qKpaTsOjGROkVY5BOyBD
81JagvULvqJYp2kLu48jtqbfGrJAwYM27AivVt26ZRelDyARFvAVu6a1nGgs2rPVHo20SKED106X
ZdyS/+7VWTXXpTb5LrjFhxySOmpNm2pEupHKTaYLcngO3FLO/keStzqUShOme3TtDlTVGslAWqA2
yEoIFEKJLCoakACIp5Kw9PUWLIgk9J0yOmezJjxoAsqmrDHaCvNX5wTlykqLBQbRUm5a9yK+P0bi
4SjhyGQ8jj0iaXvxaXYRbDosoHcuIQBiqCHqw8nq7mcA6DO0ylCSZ5ON8VRF76DAAPy/PJWyEHbM
Z+cuZrnO8PEDuBGJOlm87brZc9flfNjdNHZ6I5/ut+OSBntgL3TUi3A9C5Rwfp5t9BZ9la+HaAbf
cFpvz5CZ4aV/A6fd5CF6m9zAZYlH/o4Opaw35cBrf7qORfmFpyWLomN21/6P20kLl29ROeZw8Uie
WficcUrk5sfikufncs+SkkSEjQY47oqRbeR0gRBnyrU54coRM0UE2txuYfGkxqHlo7tm7xeI+ezI
0bC2SEzyAnEs7+iYY04nbGPig019VecTwrnxm8Hc77bxZrYjM4Ym3WxOouZfGj/ZxVLAphPsTzR6
x8Ax428l0SYT8M0hZsnuNPIFiLNjltf4wXM9y8EykLSeGRsjCmyvDDEYzlBpP8OwSKQW/zLM8DLM
iA+88fV1SxHKyu0fsxZiGim1pquLN4ZODk2xn26tVOrzLUDkWNI6QF41roBik2UbwjPnIyR+1Nxh
CtrPn+WiHsQhLlQgiq1wDqMbtjeT8B0vCLBnwWqyA7U2Bpqrsyl8ZfizkvnI2fH1DEwRFMBcWhY3
0RMCz9yy1zGI0+QtpwdFqQdAfZjGXBtXxv3u+LDIyV1YA5GMVMsuzeNlXZTMzcpjEKDqfeb3CFap
5LS4k+ldgQxaPfiCAdE4CI8H8AxSoYTDiYba+sSIv7K2eJIpoZht7PXcK2gjhp9nyD/VevUQc9hI
gBtaR8n7Ge19bd51czhl9Y+vPKhCNEe/JE25Bhw1YnBy0m1fFB/L5HJbGqhuWDF8rqPR19Fd6dXg
wNVPD82qc1ooVIuIy2yJSkRlsZZd5v7PyqsKtC77O70IGK6BuSKchK3n/epvgOU3YV/955e2J77M
o9M8Xs7g3tOuCinb6HMRL13OxdKqCa9BHaoqq/5wnJ9zwE7i3cH/+PIE3LK/doTiKUoWDEy+2hGW
7XRn5VOXb0djpvPkhiQKQfTuZGrCksjQ3bK9k4Q/6HAc6Xlp8ItSE+eWdmRtCcFCUVYFn6an/0pq
esr1v2Jw/f0IzVzkNemZTfwrqWTZTsr0X2ybAYt9T32ePDYFWmy/hcKMODfKMLYyljamPKPbvcWw
N6zVS0cmbioq7iXBXlgDSiXtb0JAh9CkS8anGrGtypgDlHmpaNpA3xJMDl3pxrJJaTOnKUIFDWQb
Uk6gY/hr/Lzn8jljEfKEddah0t5C8sLf/A9uIQzPhsBM/7kpXlnJ0btoMLuUTTDWZiJe6BUEZx5Y
VR9dpUKK8lkSczwkzwiP1SoNru3C6IiBrd9tAVvtFDTHkPpGfLDU/+9tbYw8q8uixoCnzm/p+kUr
CXJCVmLgX+Y4eWecUq9KpOAeCIaJ5nup7kHcNRufn10qmN/gJi8/pNMx7xy1qnU5rayQslrmcxt+
U1ttCwsg+bCJEWLUatX0QoBNb4i3HSjFXYFbSwK/IHdyqH65C+Zs5ZKmjwngNMNL4whmsx4kaE6T
9781h17wErrJKENX/cjOZECWTMczPUvlp4mqfdytSVgMJge2QO38Al2c83DN3xV3J1yCuciyfDcH
FCKNPjfvxtNW2c3FG8tJ4sRsluTsih3YycBs0BHwmGRc4gW1v6Ch5jluhyDUmzAxUOGOV2IJC3KV
hP+rqsT55ZFTQn1bYuIkS+KZV5oiCQRok4gz/fdrgQExb285q/xr7KlAtc3yB5qi2LuSut3QDfsG
9DXskGIp9jFWBPTM1Pw2mGcapoSPqSAeWl5yCha2yuLjRDzwdrJX/B8mohd51B6mdyXQv8+4ewwZ
kCuQgs+uKkkLrFb7Lsi53GznVPjJNU8DvTOT2p9jGRRuCvpUWJSXr0eBTX24EmiSBvLhh2LBvdF0
cruSOKXt8l5/B2mAdIaYmYKOggynFJ+vK9ebG7L5N9iNAutRPLv8I/GK1s3V8y5D7DWNalriUair
8DxCwEGxrSIrRAhB1dM0J4CxZOayoZFxslNyrwB0OvUxqW/NsVca6I+qK8Z/8EQi8+NuWSrtqF3e
8wDHjRy6V5TE41MXi9BqhaA0ttqyxyDHpja4YsgI+HVDAoy0bpV+df8X0S48V8Ph7ElxsQyTAv97
PheBsEGgwcv2d5OWE/baE0QjPhPg6cSLD9RraPuKyWmL7sAtj/6KPe5PxmAezwB8c75Dzo+MYNyM
9gIe9nFX0kjMHLvzUud8iMoOHUL0Snomik+LsWZR/bxP8eJV/6vcQb2/u9PSKf/0x74XV94zTUyn
QJ0AUg/76fsqK0nXUjz1xwj78qwR6KY9lqdFL7PvBodGzAIEtbVD6IeR9AkkSnJJtO+Nwjmm/niH
UsFjDEOMTgD3DgjshMnqj20twe7jGo0TBENvh8Evc9VwvcGVdP3hyBX6jeLg+srcCiTvDeHrkA4u
o5+MJ/puPDhVF2NmH6P//FSDLWr7MKTtF5xBr8lFMxGDh3GTxzT4T0gVHf5ZnU+cCVDULIOElQpN
aPflm7oDkRb0F4WwJu10su70Fuv62150d0lx/qFU7JNarQGqtZl9N7Yj2N/WJbXjtl34mRKJcmPi
7QaxHv+70uU3mobJwfQdPai5kc1Rg+hRqrvApSM+1MriiXNwxval4af83x4gEtn2t8qclIwkmsIr
d3WnWuOY+pip9gwA41I7Dl6C/IPj+dMQzo7TrQs4+cxDX2LYssJWdo4bKLclhEGouANTmVHkZ0YN
bUM0DBUG7A8O/h456mwDUhfWW+W24UNUUSuvNvErxo1twurWNkPvF+Bpsr+WoDM2hI+mbQhgDR4E
7D4WWuRCLikzYwIPRwkssnKnQnWXFzLx/hET0ZpajttloYOpkrS2VYPv1Pi9dlTHH37TOv1GWfCO
Hw98s8dQbD0wq6Wg4mBAw8yD7URF8ouKtbJRDEP3YvUBlslO4fY278ch5yhSFVKf8BgXljzG6J36
Wib5HPzlcHw9Es42LvS9doDj+H70jUzs5ABaAUuonUGx4WYIBewNcGDClNKDWhFTt+BcyZg//Slq
I4w/0OV85TGQMP8Z+ZDyNBHD4+7j8YE4HvlON5Gw+VzkVtQMcdR6Lkd1wBgXoU3/OAJDWQyWXDiV
eXCnF13nLKvne/GW7hb2X+z3b/hm83S+R/C8FT/EAByjf4O9WvijVPSPKVmUyLNu9a1Rg4CzWNFk
n3O//7zEmfImLJM5aqhTcrYCpZuc4dYUaJHGHKlE7WznpgHyGqId6yJsX2IJav9zQBgliueksBrL
YzsyvBxxgziXpIxDHWQUXAhNPXn9bsKNFbuR8doZ5gMuParvPTPOjYwPFhx4TVsU2H6N+UdwfuJl
DDBplDw6dq2OYnW4Hox4K5fm/9tXb9ZGdYV4iB/7ToyqJfpLQ0J2DTei10lkNdixTNRGXDP4aRLQ
eiyxNupBPhUjzFxRWc/lzDMR7ML3G9Sip19q2tJLsreLP/ix9i5i/hXDmRIP9Zd8D7vHyY+gGCCV
gNXhs2I2a6swE61fyvHPT0IVqwfcjrMoFfJBHPPv8zivMuroZEtw/UDUah0AERZOl12ldeTtspMS
MhNqus9ZgPrWBISEjoxCDpzwEtwnwUns4Pw6Ee2f222AC2w3IMfrv/tLoHQqf28TTO0XKDl5vC9/
4oOoqQnVKn77AohWhy6pcAJOdQwdxdzDLS4wnRgFOuHcPLtnLQyHpB0rtOAcia7V5G9mcpukS8A+
MeOE95QmMQ5IJy3+LqxvU2WLabUldj5E8WlxNnuZcK2IeojCpbedkRXGKSEwOCMHH5PP2EivOzvL
obaUzQf21dpGFjdfTCBfA55XCozhjb2kHiiQ8+jIiZgHSZlYll37Fu3xgQIFE+1tQpbmzOt44xBN
ilmGNkKmIfGKYKhsaEMZ0o/YcIbiS9ol1yiQj3X84mUIGBLjB+idZPfGo9C9vL8rkFhWusj0hfq7
ckgcizzxmftqPppKO8woXuBYIsG9223dmAh6rCCQlBVSkwEX0r9kdWUum5ZvGpZmTeGa2a9APoB6
/7w4V/07L3eTHom/DolCeY6yTt9sE2Tzs56J+yMIhWLA8guktK7AHDRM/DCmuoEgFJrevMoF/aAL
Ze1JfWQ4w0hWi796PwP1aIVeSGQwL0cxGgq//v5h9rbxFIqoop8T5JXDGVpyRcDGq0XREZnwizY+
G299G6CXda3tD6+l2OwiVoJ6B0HwAAo7PFyL+UlCQggAQ7dOlOvmZTGCX8zrlqdDN0ibnGiRksuk
2Yh3X2L4BN3jQBnHQXfO7G6xagW0GvEikmb5OA6uApkd6MuBqVVXcKlhPjcKT2WnG5FhA//tA5uw
xGc0JMHf2tS3A8e4DYxyg/7zHzJ70BUHms6BMY6TF464rvEJZz1YHgHwfJHyz6Djz4H06+/BFltl
tW9bbstfEthod1A6zqPMQLpKV+Aky+fQxfeOwN3qaIozLe4iR0OAatmIwF+OSspJqmW+3X8iJZx9
qWqTWQjV4666IK7EZEWRpMsT5aT19pDSDTsuF48SnpwJBCDQaTce6O5Xw5a/W8ElBHleeMld5/j8
fWslP+YA6bvxUeBMUopfheErPFqrsP5qptYn+IBJoC6WxkwSB/wMamRT4VvFsvf6bw9MlloFWExx
uqHlhaxSDAoyAYRLe8g49l3ezzpqrBwrlj4FvkKcQceD/6emznver8JZ4NkiFZUhddRRw78SfYzl
0rJ/OjsGpAbLqhbkzA8T5djEgvcQCHx5D5LjKU9AFMGBtb052icTBCiyk5AoUD/RwQFE9x9Ci1F4
LfFg4knyhjZ9MWE/pS5ccMLgN5cP1o26zjsJtU7cfLJrRmVUxiAj2Zeh8Vkh0bL3SBIQ9+YS4TWp
ii/uvr52vwB2hgSqBXLrcC0zZhFhbC7IZ5bkY6Q166otosMYyKtTz9guxdxAk7yr7hEBaEE92218
rVNwRMyzuAj8duRmwIN0Bva+7XjOZqPX+1ENPG8uLIq16QffQdhi7R+Xusjo6PG4o5hdskPkOSXd
3Ef+ARj+ghHn1+71qRmtgjWQg3V4bmG1PFRTVSKS5jFSG0fYRI7WOZEq5fxyCku8/0V5qMOyKJlL
ys29iC6HiEcAHtYFjYnZIS9hHS7h+8acHqbkYPuGKlafDvUF2QT53dtPg8to9n3eHpvv22IZ7iei
XJEWhXZv8UJk2igUc2SwCGDJObKZc4FKtNSVYc7pHKpNkO+SahiKgEhJnIgkhervILHkC+ulHjVu
S7SHGkqTQhbO4WVnUlTajkP34u2oNzAxDO7r3T6zxcdAEGlCgVaJz1qQ62N0fMHhbSjYynwQ5VJY
kWEBnp3Tfqnk2Rzj75YvFDPv2V4CUFuF7eN5xuXBYggr9jdT4rDCKxex4beyjgqJfiAa9xrcq0y/
xfb6xmLsn4pHQENP4rDeA2n7Lprdh3qxIoEs+o1Y/q3+SJnGGNYkHWStlLybHUjnQaZSxnam7qsB
BXEht44yH35j8EQmVLUKwGAiZzK7fVA3IU5UXkLSTykXA3baEhfSJWrKulS9sohO09emysL2kCGx
R6oMjWK8fZq1OeddWE3R2Ew7HQ5M+tpIPobuz4WS67KKn5sRrePCjxasTfrBz8RA5bVDXT8C914Z
bWAMgdxUN19tr/+hGgff9hqvkky8p2urkbrFwOyMuOybSLbNABJI3ifrRqV1oGw3j+SCSTSk0vtv
Edc8DxgArOKoH3FsJWA/o0EKePxzInbY3X9y2Z8jWgWfqnNHYlmnEzPJyrDOqjs5G1MtqDaBzl8n
IYtADdHIoG/WoTqHhw0oiOCILs/LSLkhgXz6q83GP1BXVqKcm7GHZEDo5B2Ejirt0M+ndtZdyRTM
aOy24JDGLJ2HaLuZ7W+awENzoubUHG6txH60SbpRn6SOXcxwSqKA3uW29O5BdPPE0jKBWQiweeIA
SpGIIo8g59b4DarcIHst6ihAKtgTOfhxD1OVyJYvTUn0pMEbQfQ56UTVG1BGr0tyxEGnrtSXtzFn
sj4u8GfojtMwwUVhIWvpiVYjcyKyryARFTDcpFco7vTdn2XhZnIan+3chANcO6m/N+eHOzufc8/8
jzkDl+p6kHsjopeG6+C4bVBshN0sBeJItig5M3pLv1Ke+fBqcmEFcvRmqA0TNK1Up/QcUzYUr+SJ
4p4GuvDfmFREytvkYvNBDpEb0WFLdbdIZCL1gW/trZ9p7vEImNT10rrm4FJxUaGHauzGXEjmiyme
lo6vRRVegqQ5lh42pKrUbaSFFC0qUECW6NpfyTw1hHwM5BJ+T6KWV6RM/YOds5de/QYRbEXkInGW
bXAkiPf8fYLMMmk+Vrwk+tk0yEe4SuiKbQC7mTFVjwzKtUJGRR20DR8kX8Ts8XAELjBi+UsrJoPJ
ssiPHn649NCJAEAjAS4c96jp4SdhxDYUVe2RTDv8+TpuSF4j0e/9LLkJZPN5DO7xbIlT1CBW4pr5
E3jD7cmfNqRXktOOu5wWfMFjKvlb+2yB2BeC/Bm7fc/gjpW/knPVyVi/h8xmR+j29s9MJ1PU+9kr
2ajzrMDaW4UmkqVfLFf2hKLBViRelZzFbJQ1wVzwJb7WLLxAzFyq8zjjA2TfvklQg0NIdopbrBqb
NeK/fLA4hLyouyHSDxQUdfYcRdAYnuzJhtg33vLaZyCtTRxnRN/7t+NOFR/NF/Rsvpl6POi79bkj
D5S4fqfXYH6BpJf0vHsSrY/mMt8Cxp5lC9hZr8EOnafNGI3I11F11WhGrIEzt7b9PJyM+0IMUFVd
EvpGFTYFp0jtCsqbAO7d2MlvPCEznWs33T8o3YtY2J+0qMe8ZIgRiX7iZEDTKhdSSQUFTBdsTnV/
Idboy7NSUmVai4mOqmJXrv93rP4W96KuqpN9fXmch9A6k0Yc/MCLf5pUJJXJTV0SH9fUegdJmZsy
unAKb0zC7iB4L6/npUqOFguSjdMKfCCasI/5dUXmL4CpeZ1djOQJ3JSGSdKqUPdh3qETVJBOMOQe
umlSA9jS7DcKRdNGruUqOYBDjHntfpVEBGv6IlFLeAefnrDnxCt9k3VWOtMp7yBMuCtN60Zy628T
FLEhzTQ0JkcZd8zA/Jwn0CDRTaYFSQOMoH+wXx7lbjlPubj9q9jHePX56qx73dtL9UvdRE9GFYbY
7gMQo6KepoT83WWjrm6Sfon0lZiubRgzNbkM53JJmfL0A7X2mWc6FWw7zfJCDqeWpsC+YSTfcukX
e+Az9l4/qR1+zLC/3jdQOu5Caoe2tTOXrv6ewbVwtMlP0cw56hR9i9MMEPthIUvQn9CN81F2dAbO
TpCJT2mHRrDVoHnxO7HH1COoO5C08s3Wy8MUnnwg2O+YM6cdBxE91G/iyGzfpIe4W/hbrd6CHp/X
ioxUMyySN+ZhP6xqMhKGDqUJQOSBXXmGt28NcIaQV2lXPMN1Zsb6hxXblONjCrnAMVw//sE5H1ff
77Ezt5XSHV3x4vEAPwA1yO3WEqDUL+T21slWjd8GrA68oedCOfDbFImHp5HENpil3Fpxg6aayyze
hnUSDapaepl5wFPUQFVot9/tKE453FPk3kC2yE7nrQkKXQZBf13lJnG4y0K2k83FdNwSvXipvnm2
fxpQlcLsJdvcCUMAyEdFp24nwTSNcnySzLYWRpLsrfw5RzpfciWpTBDIIKmd7CwCdZ2o4Ry/SR4t
BnbnZuGpnMH5EDh7mCQlrNUUVMEpd/Mlz2WA9J+Bq45jGCMqnQFB1Cy3NBmXi/mnyv1JRSZFXHPa
CkChumSOkVlv/wER7fCmhwx0hTQtZwIFHs4TP8QT5OFKo/Ou97EK9CpL/4tEnPM7w4qiXoiscLkI
qmtUW1Sc7IflLxCVOztOwtEpmzdrp5OJ7Q+CW3DFy2P0/if1JMQh9wh85Z7eKhsm55BiedAiSjov
XqDjf9y2LZ4BaeF1FLboUo/12gtYt2TYHBeGsBz9VRjyJ6T4n6FA/m95l00MQQ/FG2mwb6iWBYZo
d0ITvAaDjvgVdUo78MqX4F4hT6Wwgy76eo2kPTnYjblhRBRfaVSHh+pRQo0CyGnnqAuYkMCr/rGB
zel1Hvkj71uJCDpcXF4TK+1FKUC8U8cXhEsbhZZI62GSyKAunZcaCI+y+YmZPzLY45v68RM4YvGW
WWEEcnL/4zjLP57M0acfrEmmoX046Mnnw3h+8rtWPFa96x9ZGvetMXAXSk18HGmrxWDvte3wFmFA
xMf/WI+WhJb9TeyW5tZ1/nA0v0LGl4SNsY1OKUH83HBVoFULVSkBraY9FsYEGG5HlarbUzDIGEJ8
ZDnoGiQ8lD6P53yYZyGzhKlFsHKM+5f/+D90a36xQxtyQXOLFFhJAYwZrTbw5NofUujd8VvgT3Hf
GVUwkuuQ26k0n67hEBl0gV5EoHLNODPTwDvcbxyT0liDWHNtzvNAajnxtioa5lHycwyGsNin/Fb/
6ESjy+/OX2IYLYigoDWXLIKjUiDOMERgjrym49MXnGBmySUY6tghLH3PbHza6wSL6bIddtJb7t4r
E+TnDwKZNXweZ6hxIiMIkIsAeqA9tKQ4+sg3+/brPuHaZ7QKCmWYcnmmKFc9/Vgu7+Nwbf802HAj
21jp2ikwVVQ4wuJ3hMhxMwMOLmstECKOAtkwGsEI0cw8ISWE2ZWC2hMK6koMV4tTqdYCpVLKxBlA
1lRVTAMi8x84N+3LyPC423jCQYKf+Gq+TCMih7MvhuN/K8cOnbX58ovaioKo38frDS3XnoBQZLEV
AoJSNeUqvyc2cpNjPPZRT/OvTU8XkTMmYe8IsFyqqcUrqSd7ojJ0QfKh0evPaxScC2JbFQxnCuhE
7vyiWInKd6o2S/HjIDjhidU+XbuzIwlRodZA//pdj0DnsfYTTh3BSQRwUDHtHjPQJFc+85asNS9d
mzZnZVDqnWUcxohbumjmD1qI78uPBOEMd//0pxo0hB1gRt8ebjMt1vAor0kZDLexImFtCGyErp1Z
1n7gujce9NCJmjDg1Ghffe1OaTCI1u2ai+N/2aTGh5ZKga6WBxrD2qD/iZlxvMTlMAH6ebo9Kwoe
8PIX8oIHYKtanqrv9tMk08Ji2JDXs12w2P3t0/NewIqbF0F2xIa6sXRT3dOM3cGfw8tZSagdLwTE
3LFlinUAqAXbYE7E3IDP6MqxSkA3wLJNQBqesFGJGm+twSmo6NwPd8AVcIMjYWna0478lM0Hqt/m
YW9jZoo6ijyHKJSsyWE4Zi9TAp6xt/AUte7EOOrxc+WsoKsdm3xo/kJFo6CccGQe0pSmz2K5Ue9H
sBximlvQeIcLYW3XTMSC6NrFI84W1uEncJNaiBxcDSSZUc+94SPHupNqOEJCFuPA/tGmzPhOVOHg
EI7b7ofEZ74kAC+MayWt15zVI45yGSNPPL+VmcTQCgVFrgj7Van1MPx+JZ+VwnJJ7/JktBGK6H8F
yEsiQMYA46nkZbhJHV2PaXLLVeIQs6IwJpEjk/DRe/WJTKxg54GNw/UPoE0ao+bMbpFcXhyPXDqg
12+ja7dR8Gj04qQmTNo+rvQw5WbP+sEuYjwRJcU7VDFQFHkSQ84dlVv7UrglktL6HmJ3C2L9CVrN
iSVvyU7W0jVrp9UBe0xU44IPruQnLqm+h9vcPwoyc12B0z0Yj84PTN/PlKtCJvxzuoQXq2Cc/LZM
o765R76UmMIXEWlBb31bjnbJdmUDQcLe4iQO6f5Pztw9KKUJP10desrXv2yEEd8G0L/Br5lWU2IU
YLUEsaFliM3mvvGIiPbs0QPyjuDzT0u93PruO4ewoqCDVaRPEXWmR/eu2fqB44GWV0ljiKdWrZCv
Y4ydgBb/V6IEEnPuVptLKmyK9UNqtOKq8AYU68mJmFJg4A7MKorq0SbM0c0Qt9RfNuz51lPFakbP
KkRm8gxi6/F9F4f0dnuGqnsr8TcHns2KFY8sWd8PQQoI2Gw1s4voKu7a0KP35SYdfESiN8o814Hv
zoexSAt80BMrWpl4f0BCsoYtxlDYYbaAbmj/O492kUt52n0QfdMC02fCK9aBWiKSdDqJff4j7xv0
qepr0lE77/TLeaolFruebFVEv6FHjTQmgCbcP1P+N1Fs5569TQETOv+jQ5RcphAYESDBdS68UHtG
DDOsJGA6edAWcWBYB9sckGVkIKykXwElEcNacqAAxVQvNuPcxE3elMVZ0ijALRMHtMBP42gcovrJ
Y2JyzWjZS48SZBl/U00OCvQZ82ERQLa75skQ8yOOyCYRv3NbNA7YrySao3eSjdecQjMLX0Y4Iarg
hPdKTDzQijUnhRhPMNmMA8ejNjGKgUEb0FIRZt7k47YcW/P9q0nlCsUJsl/NsxxdYfdF+VAX/LJB
NWnIOoC4LpPAGtv5sJ2GItY8Y6+4rPYIKNjjJmX2sptDsckpLkUdqP3O8mDtyzT8PkoaSKb8Uz2o
JQ8asny2AdDyLLo4rwi6pM2jx9hgO1k+PvnJjAtPOe8fFwjThapbilc/HCdtxgSscVl0sk9wGU2L
fR3Ebxwf6nWK2HJcCo3VU51JpUlcEJ3Qb6qRRwj7CB2v1HNiJDOAN8sEzRr+8PiGRqd7md1/B4Jy
84AeiMWyTa1RJYqukC1bbMKUOvobp7Hc+tL0Q8kv/9FpLSgw1GKRM2pXCUm/BPcEqsM1hmmV7nNZ
d014vIbU1lfck8sFX5t5FhGpNFDMd70mb9ssq9zgz6lZ0JkW3VVo265UX32CvkLBt1h/G+iBty0m
r2yXF6k6jwAnKq8mEMegSskpa6iqfuqBXQ43t50rfn/yN6Kg8kdvfDkHgeAfK+SkNsAzP4HRbS7Z
XIuLaIGyC7uppGdm1MSj6lLWm9dBIoBkyKlP2KzGjoQ8f4aoGrr7+0GMzaGh2G8zTtiY7BshrHXT
vAZAasUQ68w76DuShcVeHT9wmYXbLk3CMxaIig0Gybn9Yma5/l6rXOm0yok1YAQpXsXjhLhmIq/a
4ZNdn8B37sxSiW4j5QTkDK3FRwvAT4QHAgEzOUiV3KQnX9cjDmZdq4+ZzjHsbCvvGN8OqnccEpdy
n92x13ZmBUklVIEClFsGDQen7oXL5Ae68h/q0ScUaVMDQxTPpG6QpAMuvg7UcuAQwUX9Ixjgr0e+
OnJpjZOoSr6oyyFyceDbBcOI+lk+JrEmUWDZ/z0lkzpLOSn6kpR43ZyimCYqkdxYLeF41pwLjCkt
7Khziyc9gYbHNwxZz+r+60zhgVLjTf0AnFEC4iPlG3twIORsfphSlmS3kDW3bHQqODIFa3H+K+Qy
iwCKpSxNo79Ajl8t9tqcotaAoT8TrXXXRTc2bi5MO5M5+62/6Kj2DSWt1liGEV5FwBnFeF8K2uTF
KQkbm/J3C2+Z8jPoYdNVcpyZ6NAG3CsmFY641RpfIAi6if0sCFxr+2Q9wwQ7y7VuvtTd+TvV7tYx
TI/mAcKwJ0qYDwXHMFzodBnLN95R+aWyktLYK/l8EaZBknfS9aBP4WC9VmkZ8CQNyZo69+SvgL5e
GPVPEbg88iVpTOz+NSNI47unwHR510t6k4ZZzOIs30HdEAYExrde4/zsnAGmR2LYVd41cezA10ht
QKkDOMMVLnYoxY0AJNhTYCcTsdkR2hZckJrNMMIv8kPhKVXDS6AUuHwgabrwPaPj4LLXSxTkhuMh
Ovb2WYQFBlHYTfqGZJ4QQCvK8ZbXIZkCLqIrhAp3Ldr/60lGi8zWH6ev/m2jm2a8nPDZiA34W87p
S5jdt5/LcxvlLLHDspY7hxf/Fs897ypOyBibLE9FaSqocn+lqRa7GelbvzpzipurY7IYrwAoQOPW
I9z3558ZEU+HerXSbDNeWC61p7BBmEDhvrXxg5MxC0LpaN+N2sfbBM3G7fxcX+P4E2QStOFF4WLU
UQGj3Ux8nmxj4x0NjHHNGrHSlvq+HlchxWAY1wBamYZtbBAEK2h8UkWqvEPqerixkS26Sk1v53/T
3Dg8AVHR2vhVJKMS8ZXHD+VNmqihYbYI6w+V9leLTrEe1nKTfZs7muGOncxOzO8JBg++tMLWa2eq
AFNkpJ8ff43DZhmi4MN72NZok6tZmzCW+5ZiNRK8G9neoCjyXjOTYCr1ZVz87k3k3LibQp1IU4Km
JppNV47D9+TnOBGfP7lLVAcOTn/KFiMWFZsMBBFJV10ExILEe6dsmitm+0N5US2RenB1PYopOuB4
v/vaCoFCCe0L88BQQZWR/3X/fjk//xQb14TWdrkDmGgRjx6Nlm/O2KrLor+bx3ysJM14VcMrw6B8
4Il0izpRoGqp5fPQs0rdCfIMeXNT4rvg7dlMRPAfdTrOUAQ7LycVzBt9sJhTZfSsJiJzuUb3XtlP
RnWAPdq1qiNnSmL2a5NznOfzT1WbYCPY62nxanNuj7qak9eFXjCr1s7WlOXr8dOLSlCcbYtQfr4u
MDofgcrfFeq8Jz9TGhX7oVbc0dFqOXQ6+hAVQEn7Hj/qAXmww+xEonknBVTkaIRcDyJKxwzMj5tA
4mJivJ3JDcgkdkcyT6uIG6XIXylYudv3zV2AynL6EgFoOeMGIaEM2IssQKevxlIlPSgjejtTOdAC
DZCd+REGuNBk2aYgQYMSCGCpSTZZwFA4/eD57GIirDuR4+zROFJw3hAXGC+HyzkW08pgO5+vvqDm
eBTqYs8DkJukmpWFOu1qmm2yQ/UkMrxDZeawz0HuCI1X/t6mgqu5r7Zx50FTtrRr4aJ5UyQ+Xljv
O0CW/12Hup4oJdi05JfzE1EL6w3EzEMZ5mITjfvQN7u8uwn4sJ7uxUGj3blgpNJ6HQZKHS5LCkwW
JTaL64W6aS8P4FovOjw1sBV/uQWzRISPF/Oku4RlR+Eq+nxV9zMJT8Sa8PysdYG+DcYqVMBHucHH
nyEV4Rzv8HbQltsnKwYwYOkambO73QNZBsm1B8rMmwvMwxwl6DgQSd5ADF8KVtOQbs+8KLhvKgHE
6XJ1hx3c+xmTaSeEcRB73j08cLdGQ3BCIgkQoM+/uWhUlpYtxbEawiVEOnrBenI4/DyA29NSXIEZ
8nVlrDbTmoz0gGRcKywiWWgxbjiIZqB/VgrP5MNS+05iOvBL7V4dLGixxEqM/sJ2ZSplIpm/1ZkP
Xn+vb6HqXcuBEd31YikP8+aCu9MyK7Tv8WGi7jR3P5S8H8AofKvsDyzwtbrajZi+uqVoZbFd8tuZ
nZ1kk0hI9za1avyz9kVg2K6aVuVWd91hxRyNmlnRWlY3HKrmViZopUUgxeWYbSBj8AkXOxyq3V29
mNgbFGNc/A9n/sCdfAqSNy53wDpGGP7jpe1Lpgm0+OAeO1Oyt7U78IZpN1aoOsf0WlZKsL6+Jy4Y
ZSUu+PwxSgUtDFXeNlGFR4IqqdmLc5qNWVA+HTaN3j8Jao3duqxjKhAwnjA5Ze6r3li13cJeTw5H
GN32wKIzrDDk9rFI4Xbvnjifxx+niFShFxZ1L9d5Nx1CJMy6kmLXmchFDTLlVJ7h0/GkKJDQULsV
v9Bx9r0nxLPH8EXJiK/OJMqwtAYNLUAfoDUen7PqJq1lFpRVjt8fRXRf1zToPKWlwGs/TvRcyamE
kKNi7bsSz+EaI4XWyu433AeZEzVBnY0WEk8AqiUkY7i3ibWo4MPAndwI3EwSsEdx6fd1HwdK3EdQ
Rzw59I9q35EJxG/YxCqNof4KTgltG65I4FE0xXJfa/GscYQqoPnOEASOG9bRa95Zda4po81HpLxn
7es/yXN4CzbShRi3j6Ng8uVJdDZ9UCzGPfZmq3p+vRtoY9ItAbVB64XB+FYbod48zAk3lxu6XXsb
fGVMK55VaUJKmoZ6/gqiE1wqbsu1nvmgfeXqh+61Bp3qwac+lQq9OxxQ67/g0kpaSs3SCxSctvY2
cvuX9zM2CgaAWmPi6AM29x4jxrNp7Iw9NnJR7IBWUcDORarMGH18iBSV61mps5D7GmDopl4lCyor
Xxp1Q5yOrMWvWwS3e+iw6RieQ755h9ZbrFVP0Qhi49CqsTTGOUpLTatFG9fabbf39fBc1KeTzY47
I7yZ4DrYrXeGea4kyTVKJt+pT7I/S8EvuSaNeJlx+8qlYV9AhuLakrPVeYF5d/t900JvDmGmcBQB
PWslaeNOKdJlG2RzhQxT6g4v8iFLaMk4nzD/91sLKR5q3ZRgmkOm7+zT+S5cfMPUOF6DVc7n3L29
42tLStzndF05gfO9yEMOE5LBm5MOLl048+Kxf2AdmtF4rhPAC4P2PWvtE4KLsnEHIyRK0LJaiJW5
FlqxPPklPfSXgay8SffGxgvcRfNIQkhauNFFbB60XaqexG6pIlShIeRV2R2uo9oM4qb3MtnjOStG
yf3M+NZp+ehXZF+UkZSi6CdaERgOc8qlPX3pjjt1tKG/eHtrnOkF+NMVbz4z51S75JU+B53GaHB3
GSDOxJVPCvIO/iP0Lp6+jcvKhrYvjKAhsQ5EDUAvNwBhVjyOztjqmXF8FwXEDG05KkCDoc0aolAa
AOmY8xPsM9UdQ6ft8pBRXXecaSaVeQ3399sO6wYru3IupXoDN7UXgSI+AjMJ2mBC1/XsxIN9IAUO
9Z6lDW8Nscb1aN1IEwoVoW/4ct36QAGIQLob6N+Ky1CbRF1+0/ug0II3jLVNu9BilyN/eHF2LEIM
iGRhOGlvT2lt+rtjsq5fNY2fEe1X6ZmOX3kgTAOBsM4tnhq4+aPr+v1KVr/gLuzLz2SgcLeLuDJY
+iGYSmaliCbrXt0yjRPYeZCiUIMjCYWa49TasBA9eT3J4cLywc1ad1IZpv0qFF6wt83UBkCYx9vw
Y09sLFSdLU/01gMTQw8oV02BczDbN2NBX76M9u8AeXAgQRh/YXh2y+8lPNH96WXLGUlwSPPSWmPK
uyacDshsgm8jzXoUQvenn0VIgrGXtXd6qT+SIIcC1QNnBXZAWE+0SuNMw1AMqPznNXMePzt0radv
PJ8bCPw5vp4UyELuQ/na/rWRILiYCnF2cY9uLd8HOYd/bPEjAfSKkcK3xs4m7XsAFEzwvbZZ+kEm
AUZFJvNccqcEfh5yQAovXA8QFFz9kc+m+NCBIHR0n1rp9dW1pkfW5aGp5nFbV9qkzYDf+gacpWyE
d2uXzTg1MetrLwFOt6kbUetwMEo99ES6A4YpdG0f+fC929WH2HkeL4FyJ3FHAwUu98U0IgwDKEgx
m8vV6LOSgST1Wed4+ERPzWGxpxTF/lH+ITDYleqW6HTDNdB6k8ua3Nth98FAjqDUEXBPiqTt9n3M
YUUHLKyRe8ImWBHLi8iaFWaYPWp6dnNvCQ0GK67tCoxX5qLdxW3V0LKFGEC8TxZFPFA8e6vd2uPp
mTaf9mv0vck3oS7TNgr855/P/YYhU78awcOZyrQaCdl30m1SYYbE6JtbDiMlSG1ENFgO+Q1MwbFp
FxN9XFc0xfDTMgBIsy88dMQdWiEw9CnTR3PZ7GxoGDyxGscmf9Im6/Xd+XMYzuJr7Yho3Ce1FtGb
UHnxXyLn9eWB0GX1UYIgH4IMsS2Foa7QdoyHnEVdwzYewiZ2y14BgCuZlARJhWxUbX1winpi0Ogf
3zsncFcJaEQ+t7OdzlwMus4kLs1drPeTiI7JMOY2mbkK6dTbR9UcVty4lJ/lUXLENxj/VhOARqCv
7NCO5Aibr5YatdOzNpnOBs8lc14VNj0B+F1aimpxjYi8Av/DKvWWi7LNpjvlkWlAKqVjNA2cSfsC
H/XuKiPYQ/eNv3SKJe5PWDR+gnPXIaMnhP3XRaXZ5N+R3fNH4mg+X5tbuvlIsVQHnKY2cnNhWmg1
4OjY8j/twbWqHAYPGebe8F3l5rr9D6Bns1woR3t33k1pvT5QyFyyjAhzhZ+c4QwKFSnFM3RaaWPo
X7J9Xsaw2O0xxYCiYxCgeLQ6Be0CjPBQbpA8zqmQOWU9PncBA29UN1HqMTY+r/5s/Kvcmk2pMnUb
PwQaPx/UKj3RURiS9w+u2Y9vU639aLsgU1+aDqvN2FVbD1RGZPghB+iiRoeI+L+bngv1JTBfMElT
SUq+YCLO9yfdyb8eVr4uBEH6HyUFhSZa2wtYLzhNplIfQ1hOQ47C4ak5rjvP9Gsnr/IQhcJe8sJd
CZ6xMVMDFZLVrb03MbpSZbJUdX65Ui2Q7NmOldEmko1poOsrR2Dd2jY6XKqgcZ/06i3rM6Bav/L6
dLeeeDsoBgCSgo58oPMYGJzKTcwbMxbnzrYzVgzxDb0Okrv3mc1WwwxlFQjaVSjbuSpOwE0Jja8m
BWH16RD73nyOB4M7rdN1OJzBxnt0HIJREIi0SPkV57p2E6HsOEVM3+HNqIXtMtjV1hZJNgOp1VO2
jtKIgGboaS6d4Qrz0SiJQaF+T2OVYIQAIokwXuZfC2PooxB5IabxKg66BZafFDm/NUYWP6jIkwol
VyFjAzbWiVIZdmJfE2RqjZ9yRLDtaAM8l3ZVO8J+DpogHe1OTaMxuVsp60WuBi6gqFJtQPsY8Nsm
kg/fIGWLViz8H20DeyMe1EdAj7ZxhJKsaCzwRfO/5+0MWhFhSKGf4a5N75+ji69cItWza5FT0Mqa
AXhwwYldmvF2RIlR44R3XKOiNqYM1a0uw3VdG8wF00vrAhBZYuD4oLMSn/WJ4yeVdewQ1LMMI5sY
unoLuA/h2+1v0CnW9F0MCOCK9Jwndl9TiayGHSq4s2/DtnPE0lKdxJI7C1XSyFUYvv7TwE7QuFNY
/xvhZoBK/0xUr2EEfJNRiNXOAPNrfmjrKhq0K1NB2BnXcBPRQe3d5L3bvHxj8K1HyJ+HPyKlE3CS
067UZH429jUgEcrKnGVFEiPwxRqaHy+9fB7sa5EKN9Ge6q19IZBCia+spIa653D8VSWD8H4Lo9E+
pk1FQANz9o/wCkhMhnMFxGOO03YGUg/w9bjZS2Yo4dSh7VwrtNVMFQlomMJSDT51Z+woeVCKBbg1
67QZ53CgJ++0GVWuznu+RVwyrYSxfuoPngWutekeBi2S2eU/q6uoriBUkxfv9kz8MgabnHQdYomA
PsvKqazhGdtCAskMeAVk8uWOyf7+q37+bfH/EiK86p9SuhpTcwRcvVby7CZQGvC+qRQKrYzvjbIx
pR1ecPFx4tAER545HAhl9es9gJVJtcjGwRL1hT06c3tG8/D/KDzOU9rZdo6d0orFSUq4NWo3JG/S
IoM3FXeQb0ickMQ2oB0WddSR30g5F50oasP+rXNhzyH3shJBZuNOE+e5Zo/72c9cVMxI2LkGNitE
yX7L5M2qBFNinGNiKohWKPBzVChBnwJWxjPsQqp8gUnq/uSZpnAXPTBJLhWeYK4dMFfV4G2XTxPF
4B7cQGH0A0L7sFL0w/CsUD2uw0+jq3C/CY1TtuEODAzMQ6eDg7oMXIWoW1G5PqI/ciNuyHHPyIur
xVnoSmYvxCz4GWIht3Iau7yvigz0iI7z+zjULpJVxclJEym+xrhgbEXW5XJeYFHvcFdA/DOXf1NJ
22cyCX5pqhAQqW0oDkWorj4nKv1HrXdWxSTLSFKq8/eunOX2PMBS/NLbbnyyfDiEKdapbNa6Klvp
GeQSumfoYV0Ow6j0MPCOHGsZaei9mEzNEmnnPFUlVYO6ZHAOIWjCc4aOWw0trCoY/sfOj0i6fxdd
AG7dJiAJRneWtsF25cI0OMcjHWo2CAfruqktiM+SenEM9jN+ClNW+c0SfuBBgSd9xe1QP9xLnHWV
yS7c8BRGaj1BVFfhW7WjLY/AwlpKxuS6+b6OSJTr5MQdRdqStjR9DZyuaLRTjUo6f/iTKhEeSjo/
phreFmBz8qeyf2H2IXQg8IHPTSQtNNiC8P0LL5MMz6cNFMMNhauUSUN2+ciYJwBfKLuhCOYyA73J
3Vp/PUiwM83Cu3stszYm2KD67x2fsZuRjTJyVpl84hN6CViwkiL12UiuMPMHACbb89ky0cc2szMu
B7joELYcgdY6zgqX1KxNlsGCqQv8RuapBzj8T9WtPSud315ofgWq/3XMSGXVbEIO3uKqzW+/if2d
WUMU8pHo9BqoVYhIS9zGwKEGtOiE/Sacq9JsKk2LvBtw2ppzRGtgOyvDoXVXWZIPUxb24TZKkKyX
8s9CJH0zm80roaumRX5Q66FftO+rHoGtEyqPKHQuoUUSEBP1CHGT35f8W8JTf3WX6QO3UElYbw0N
0eT4o8cmznRSrmlgL2uHve5HC7MPMkHnKUcAq9+yTuucr8PCSkBKz1wk4SubKOk4mm6WEFj/l2YS
jv3agnKZtKGAcatorSp9HeWyKmLScMM0wXFY9huNU0L1CztG2a1K2RDIhFLYgY9T70LBVV/wY7hV
lYGSRmKetMR9i8O2bGyQM010zVjIdtRFeidb4MWjILE4a2zbXSp5NqSF3BddW30k449/HeaKtvd6
MOKpjczzcWg3GFoD4AacWQaMf+GncjjwK5QBNdIn908pDGLO5+HlNCyzjf0K/T+vRWxzd2Vx/59q
0zJZtqglIIWUdMicx3iyb8Ct0N+m+x6GCC/GKJercOZxsVALrM9QeuWASSkIl/ZwBLOvKfPjYjgF
dvRGWZN64OMQoAlxZFMYmCCh1CVPF9+9EVnHAaWglItWLgvRJIcQjsQwOCH/tZpqNl+HmEbfvZtG
0932mrJZ4yJHXlUq5soy7FFn17pglpUe636FrEketCYvOVsadjYi4TwOFJ4iIK6QViBT7rtJUv/D
j6Vvx4RQj6xVBrv4Xb8rIMzQ/fcCwi2AjTfhmm3GhzbMfdoVSd3P/Eym+BUjn+qVKp+Sn4cpEIYw
6bv3aUiQRu49TjpdgKqv+d2YcgnrEvmoBYn0Yh4TUeYoglP7TPoAd05b6H7oe/ZuYGUxv2IppxRW
wufhDy6dJCY/pX3HBYImDxzdrUNVuU5GpGAJCmFxQNzxjHBD9geUsWYSvEk/n3r6k4nBQGN4rCGf
yBD70+yWEFI6mjNFnpEs1NX6AzbKbGs21gHzo4mfOPpHZ7aPxF/o5ox2NEEP1TyEqDVfPYLIpFqJ
+oPXwoh7anlTOLKVTLeLl1s8pLR7zKfCBm3DRVOYtAFDy5IwzjUL4IZ3ia0IGYU03acYn0qVvhd3
0+cVzi1nE7wdSJH2seBBmUCvj03XYDpoSNGRUuEWnOwLYc15oYilOP/LhIFvf1zGyC0dFMKezIFL
cg4kXLFMuRdB+oqgqsAy0tjV493RL8TUrCwB41T9zSYDkeM9OHphcQC/4cZA3KOANjWzimlci74S
luPlOWfBGAwBuRhu66LLvAuV74AjmAtU6GwJStm3KdkKN+x8PwkL9ENRZHf2spW+es3b8sNM+IeY
bKZZOAv6RZJx9Nc/2MqpWjdJa7GRnnrf/pvgfd9EEyrLhERQ5dupZNqc/y8tCW8gj6YV08+y8vx2
ewoT44ejI/CF+v/lnKSUA6ALhtzTog9Z5ey/WaNJ4f0HFGwAz/ybzLUmP/u6bMD01cbjmWjjD/Vi
rMstMvo8zvwhpvT8d3JpRCJkmxBcsXkq3iSaIipt1e//Qmp+O8LEJxICA8H96yPRwuOLRe9ZCok9
844jt6p0ZvqpUq7S7HjKhA4LATULN3Qw6u+/r02yMB+zNgXfB/OlnYcmtNk6ae68bGyHtSpaHsnT
jBSohBrA/VXAncuY+RIe4gaisX5xixtbtzZQFcyl350zMEP1sICfk8FHCTRIHMjEfDn6B/gPVhMu
AwhgBvL9l0uYrMAWGL85PtD43PqbmPcEYTamRaoE5K9qHDEjPv7H/SXESE30wvpsjl1uOQzUkjEJ
aQ5PTp9jjfa78rSEV/m43I37uYzDhMrqn68pFJ2NdWydl7DlZTvJveOuGw0ck+ZGzCKV/l6JzKt0
V6tDAG5MqZdO275sUWh6hWlVuJ8BrOGGF3r2X1A6a8Uo1slZxE+dmT2EjcbHdej7F2emSmWlOWhL
zYtwxS7hJa1RJeKC7rvX0hGyGlpStJq1d8cJXHIlZ1i2JD2VIlLCsSES88kvvS1ZC2rXSVsJLFVw
7Ik2+Dcj1gfivQ8DNnqH7zT/QXTYXt+IE/U7sSCffKxZ9agaric7JJvTKaJdGm1cdQxQOp/CvVof
tGNlBbX/INgsrASUM+t0hVzp1bdvof2fRasEaxAPMCOYoTD4v3T19H/w529NzjsVlB7Iit0ixirH
XJKsS5Uyp5hsAFCoGVNhsImZvS/QZA97duDRDy8ijrp7IC9JXyi99j9CqzZ6Crl9UvSh20QJCt37
+uSYABa2jn8EuzuoDhgpftIyx+FyyUAVork3++gdFwp2wMueYSonWGEPLUrz3KPOGIicHhT1Ue60
OvQRqomo6bqaznVTXkl7Q7MwUwwYj5zMgcveUkMvv7xglad8p33u5Q3UqoreFnr5wl6wa/AcvB4x
TzZGpFB90qjpvWycwxD+hOpLNlAmEogTyP4W1VlaUChLB//Yg3qKZLsoOMWp4IGFigt7buAg+6GE
yvDbuGy1weB3lC/vTnXFRtG+LOxSdQhVDArF9F8RUUvel/ndqimdCLldBV6/fVk5MJMQrKAxjhBA
kvOnf66enP8RkPDCIRh0OO7XvopUHsLaAg8IckzojcgNYTO3hkNl7h7EB/N1sdXNOB4alnce+5mW
pw1eTDFJ1MJzSHR+UGF5jUruaFvqJ6UcQpqsUtJvz7o7UYvlJOLKQndy7u/Rr5BX6Fev4VHb+93v
7Hr6uJkoc0z7y2lXqVyKQ7CP54F5TnYyPdr1ysO647rzYtJ0Eby8toLWFWpQf1MpqGy8FLx3UuK+
e2msJ224+eC2hup1HF52OZTaUPhsxgwuF4iEfhmjIYd8wwrXUz8JsPtrnoHLV4rUm+TCwAgBvUtW
qMCMnTS7de40GKonGhqNBtEJPhgbz+1Ebh4p6qz3lOSXb1jEWenXDCVQNKgCU+VHDpyzTO/QEjVD
wdzkYWASQc6hwW5XuieMgiHRBXTWb1ncFcqqrQZDGQXD3CQd4o9cl5/DZe/a4VJeFMJaZnt2HPh8
l2sIhx9f0yKMG6y8jCK86jaWZlYhYBea/di2K1I7HvMSvfoegakNT8NtTnhbWQ+0s2gT18mFpz56
lPhITtVe7fDXX4/3B/zyPSaH3SIAbovdsHaOurcom2rNi2SUh0vNPxPuOFwDxFmi/9//8Y9BWFkb
9jmMI2w0cTSCzORS44R0mmu96zuBzpnBntMagIBg8Wt9HclFUJe99cVFckjLvhmb7Wn6JGuXOqfN
PBnVK/9RIT35wlQK1HN1UrYPkMAINH3nFkB+s5DkbjNA7FjZ9/U9PzqaVmT6JWjdY18nQFqPWDrw
ydHRps5HrezTyJimCQ84hyriPLnK84ILcN8c/yi31jzKHeGTTBl/DCcf2Tct1+GISgvo0PBztSwq
pruq231nzv9Zxo1S8S1IgBbODDoCWoHdKDIxWMJuB9IfsFm0i+7zyTffIDBa0+TuVjuCa/+jtpGT
MfVFLgGWR03ZEn+CKQy8AO2PjnxtrbM50QsTGiMzHlCp4c2GUoohL+XiBgGhgLji0ERcpI2Tbynk
vVUeNG/b7nTvgrYqUNyl108aZj9dfjHILSqmec1Mqaxh9an11AbHF5xo5+pxVhC/BAEMDScok33T
y8CUdAcikxXcS6ZNfWGLBvZ0qoI50rmS1zDK08R3IjyYWSZdWO/s+VNqcB+YcKhzIHnCWz9c3Fnm
LvlOa0OkYzcxqKAYa3xF4IjWGHtVpBCqDIHLAtDBaBkcaAxpOrocYoZ4WC9Cfm1WBQT+jyNp7HN6
neBWHOkcssbF28JsKB75fQ0gJekLRrAmABH2tIuG2B72xBGVPk9Yldjeju7p7aNNYfhCBF6tioJg
/dM7yrn3bJXpSXfcesqf9Q6rua12okrKkTN0wnfhY5dgZ9RYqCn6Vcay/eejBcAodWM0YJ2BBRLe
nm31TYUFwSimT7DqKb/gY+fyO11DSFH/b+I/gzKDolBsWX+RIM34v/wQSwT7Guawogv7YRncE1NG
N1f3Lsh9pibs+XPK3C5yVOzM4bMI0fexT7QqSFDZ9r6+PqfU9JirZoju2NMGLgYZ42IJpSbSCEQO
VZLbmgki7ov7W016K+BZLZ5TUiTLuI/lb47vdwIVUgUUmP+9U5+cH0tEvNHgFU5Bf+QF9NgBKGtF
oowO5ECu2pcpEKyaQDqDJ7Tp9dhUi7arrHRQpDNsZNgd43cS93gid013HXXoi7H+WM1c4ho/m99a
qrEijCze20d+a5SNaWXMzk5vCzbY/VIv9Q0itAmGg0YJIQ+Z1eRoFeKX8bpvctyjyswp1GDq/GfB
JVvwopw0MrDu9TAnrInQ70qZS0W4DUNbFJEpiNAhU1dm4Tf7v4Wy0Dp73cNDZoD13U1POnfTBDb5
edQ23ErwzTbh+Kj2Xyt3BMFpQFELc7L29fGlkrOyhckN3cdHG5p8MzLZPNIojBkwd4xnnl8y2A+0
FHM0EeAwn3J51e3KYChvlH8SQkGJfO0wz9zlbQyUDFd02AURrgVuAYRFbwiJLBIfc6t7xB0Y50J4
bNVQnVQtWg55/YKEKIeWktn1efWg+Eho3PfgbUj9xL20KUJmtJgt7/rYdVGRatWbij1Iww5NMQyO
qKe+xi6GpBJ/Gmh5OtO4hCc219jZmf7mr6tsMGPRzb/izIe/Hf/EdtohvNwKt9a/vpcXNoV8OXiQ
yjFzVMFnTo13VYX7SN40SFc/H8yCgPnSfjp2slaDjQ/halGZ0EpGi5Qo7Vr5GkittaSFtfkxvbqG
HC3nGSXN8gjey7QqDDTNgQPkXG50EP7VCKR3xSdgXBShmwe9tiGElJOwezBnE7tyoPQOqyOYAZuK
WwbCXgl6oBrQJ9zFE8elFRankiYRkuUl+8Ky/2Mdw/rC53J0ZSTHzHpVFiECAyoDcsZfz/OTEict
vsMmsXJHROBh10OcNRUmlxrZL7u9TC8D2Zd8SLjUPfYD4I57EmZ2n5yibL+BqNbpYcnZPT5Q/bPW
BUL6aEHVfp9TUV/79sdEPZbOFusN37tYH5/+nNJakVWzZO9tNwcmbdNTv+kGPFwukq2yoTMSvAvE
LnJrTfnT+VmyPvb11i1ryluoxfMl0gaigldEilFEDK1Aa7CQSQuUsJtHKH0QrpO32wU98a2Rm1Av
z7dylR28mjhZ780F2TMCpTDxqdSE3BkGf8L4D3C+mWeLlSTwijHB+Qk9GID1nYIPQeAmutMVq3T8
tH/pqD8Eotz0tGPEbpx2piZfgZBH80P83siHeGAVmH1J/tSX64PIWRdZjTz3l++7vrPqe4bs6lXm
3gD1LbUgwJtaRea2m18UgBjmOqbUnWLa6BwJxFQkbEN396rpeMXw3ilsoQcEcuqiJYiH97zUylvH
NroTmf9gga5FVWrkqDYSyVogm+7aKUFainhQWO8n7TvP23P1kyTuixvPNaMTxNXflxhwuQV5/ZSw
ZymTUN+ZlsZa5bRfgZYsN2Ej/lYe7Xy+9ud5ETcGagpoz8kLDQogPBgMGnS29RvU7zrC9cmIQHVM
5O7lBWebxXGq73JpM7jsU57vwo3RxE55645SJax3uGs1ijs7p/57M8LSCVuUOkepaaSGNIhBOGJZ
XyFcndv3UL1BkePEh3aYdIin9AHhhIQXrViMYvtY62iMEnZiVRxdCJp4S+H5utt5lqlixmnyBoE6
/96WITCwE4uX2VGyT+6hExasmvPxb5HLl9G60rxEuwiqrK7BMnPKDNPxXh06Vz53nsVCoJ0CSHr6
QAGHBz4AzvuqA30qDctaBfbfJR/poo55DQGX3fx6x7ZIayvQbhVyYPeuaNpeAbEXJW6obdMBTwTl
NgkMRcS7CicATtHaBjTVX1nJlM782B1i2qU4QWQkeYm+1YuHE3OfEjQU6NHFnfkQmyQImGwNi7XH
l1qKLdO6XlssiOo8YvKWkNaf376XY3ZKEAHx3aO4vxFkqq1obEg2vbakyK2xrYZyjag1w0uIj95w
teT5fG7ZpHa9oM8Rmdr/PusOPEIhdE/u48GcByhAlQIgWhs7ijSXIOFgWuIpU05qJyxs0Nwhig6c
TARSz26vRfzWjzsKXhqKsI1sBAsdn6gWzWfcKgdwxzd5N/XBXDjIZcG2FrTPWYKctsWYzBPvKxco
v+Kl1wQxh8Clx/WChX5Orx1wzPplVAlU0i0JPgz6XLe24a6KU700jRghyDSZvhL5erUeHz6guJ+r
t770WCUH+COhYsVQE97v5+MHDf3XOyg2oMan5TDsvB8RbUBDa4eKh0oBWZSKcyiCEmYSdVUgXxSz
smefA2IQhqyOlMfD+IoffNGRo0dyfT6a+yrv2IADnG+nyd1AekdBKBa/SzIPnfGcmZosrlRyCpBm
1cfRFV1Kq/5+i/uihs9Z4wkkBN7YOSebm3ejqzSboyHKzq7SWe+nSteYMFYKwRSLwRguIilHw+z+
UVdyBidfIZQp7DIcHiqaCFsytrsvftvR5/Za9c4UR8kwxK/WIaVIFj17EgUHIrwZZODkWUBwcwYB
qTgpxz5szvIy+7YGEOjJrVuYNIyecvfScbmg7n/dHJvOZSCTY0db1COomdp6pCEavmVfXvcDZ8ga
O/ARDMNnIk0dHuiLRMHYYtCYacQd1bvH7dAMbplpkGye7Cs3Oj24Tz5NVw+dlHopyYX4N2NeqD8F
jW5eJ9y1sN8a/utEohzJvp+Xx8JkchUxh661bkf7UOTosxtpqBFRpVMqpLjP5+SbBo8XAiUg2xLG
v8VM/E/7YfQ3waVQZFoV2P6NavCOQSkpPtj0fa9Ta6oIFeiFcronCNyw0BF/8I1A9WTSCR3k7Fmy
3ku67rmdamT18Pkw5dpCpjN/l5mULjfaKUbzKeD21wXwNawIPZMaRqjm8XYVkHnxI70G2l/kn+0K
O8Y3lOkwoxM/Hx/VpDfRz7tNPmSkF6t44xrJDV9ADHYF2M+3hSe4WqGb9xPG4gWHnOwCPSTOdQuj
/Fn74Ggmb1jYvfuVGPiwk/ZM0tsF4o9Lxl75UzDit7wth0C8WPVIF6roYnb+HoObYdoxZp9fZYRf
EthhyGhFVfHlx9UE58ZQpwL6xlGHv60GWcyiCqBVawanCEZp/LaIG0IYZ0DhBzB4FYNdk57xIS4/
t5ceXSKDUIJ5Prtn5hFyENAtllTgM6kp0ZZMiPCAHLV1Uzhya8t4KbKN9b8RiSilaw5uRfSS7JMS
rvGqUTOMkwsENjBZl+ODGrMNKCwYeHeUmcUjJHMZqPagxsVDHQ189GUkntTp+ym+Jup8HefB3uHr
KFXxC8HID45G9mSxOLYx6yY7osA8BVVRzNUYhIxeSZlyP+MfOODW8BZNKJdFF11NSJ8GRTnpsao4
DzdOjKW/7EN/F31gFQodmb2pP0vS2k30if8Nftwz6ceGT9KCcpzJuQD/KnW1Q3SdiQntigRBvtqS
xB55jhWzWxf77Dmd2hU2SHlw3iUlZM1tQEuAES11wUrhZmNzgZ/Jcs+g18ubNo3dGLS5sZviYSRf
Oi7EagWdU2eNDXXtq9aGPEutxULlDIrGLa6TD9u5eYCcvJAzzciWGq527Ke5fybkUKNwRoOGJ7KY
aVJtAhW6OawaziStpf9DcEFLdHFOPIRWcW9lWSuSEiZL1UzcDJHCDN/a1Nl0Oyfzn1Im1GLjdgDj
lfZdQTNYarY5Eu1AB24+lBN95L+7MszNV0fNdvRHw7G86qODA+78yCCIRgMP2TeLbzcBqJDjMrc4
cXah9y49Rka/eJBpC/WzuUTzAuc/dKMaK1lPmO77IBOmahjuhM1f4U8W7pnhaa1YPyjKv8FXKtul
bE8NEU5VFIaEMM7/142dOrA+LcTj3nlX2u6qFuZHwYnqLd0pTq7ebb209wKDuS4PRk+GU2JY4BKQ
u37JpPbvHzmNWV9Fg/4l9wOw3i+SnzF1BDhQQ0N8cigV/57iv5GtVqK4nrZ6hbj32aAcPQOYPxNV
+5IrQMH52dePTUJFocPwO7mDa4nNuHpNPYzJ+jO5lFy+i3Dyf4LVQRNDKKUboFLDOTJ22M7Wa4Ph
YJh9FjW3vWsDqu83ZEbFaOsL6DfuClyCqDj5mUvYqfsh+ggFOgBcJUldTX3/7Gb5enjmfSe8SRbs
yNj1YVDmV+jKkEBg4fC0WEX1pQv5sBhT0B2Km52OA3WBJ3/7tgnttbsHpb3ZrzX+CLUTxzACbKSK
PwfRnB2HDu4FF3JeOw5uYPvAy7WqFVLVxeqX8I32cAEpDIGO8D1Yt8IJhGt25wAIn90weYv/qd23
BiYKeBQ0YM6w/pKZD3YeS8wKSIsZcC+bsNOouWpb6rs5ZkGrWpb1PN6xXpRpBkycTeqU9uGCCoJn
ZgQw9fJYk+9vP3DXdmwvDDnyOT3aERnDbJB8j62mhHjkFXXdgHlDuK19cICBWTg09RnIqSXTH+XA
Y1z2Yb2+6k5BQKzfqS3+nHvdtvZUx9bmh1mlckXsJuWg0Az7oxgR67/wiBRe+twUbAq/h+N3A3wM
R8Zn/g3tBJvopqDDHVxquzB92dZ9W5xAfMBUMWa8egeK4K/62/2Cj3ONQK//e0Or/oL/97RmqMhW
g7LNOt+JPYwn73SvADocFV5sgdkdpwOZNW2lWrqDPNtk1HQZn3dSA7ChqzpMVZ3NiAaHUS8/iVVd
iWYEWiMQLrJNo4ZluaZhVLfD2WJ6BX6xmdNPiB2VLynwwl+yxIRMZetmOt09YSI4scmpcov6jIrJ
gMxR+CEcOCl9xIpl+FTZhqmd9ctgiC6fOfiCZARchLGbb2aWD/RiM3IsEo+jWugfXh59BeDTgJ+y
Qh0gKF2nSsSJcnegaMnyBAYHuiaPC9HL/6XHp5/9lkkAvavVnJrbnwl3a7RhIMfc5KOuZxgQ0ls0
9rJezvOKu96BNmYUIo0e1t7gO4rMdBa12HucjJ34tDhJsiVMitv49AR95MVe/ZTEKiyQKWZGoTJ7
a3nplwcYO+r1nmWko9/Q7PuTgVjHOIvxo5CIqj0BzVvlE/409tlBo49tTbK1LXt6HU7b257bIe3t
2tkAoskEfdA6H96RHj8KGLxPlRFZfVjxaII0Q1kZyRklhJ+PLQtRrXI2+WKZ+cB4S87/0m4ivc9F
tSldbucnFx4nHw2evgC1aHAUTf8UzzzaWl+UfAbX6Vo/9YmKpW0uxwmaEWowTCgy/DUgFiKFNw0n
gK6tAewvHartlArzexhIOacmPGzWnu8BroTBip0jbavDKrmLcaEIyPoSKy2FtybAMxyhIho+CdIz
QAJ8wOJGq7BbFsvMQVzMNywd3lh/uKMr7jYKYUbcIBxzb2NgjwksI8PS1xrG6sQk5BtJpSg5K5Rk
tmD/hkJF/CfBfzaRThVZBO0U7R6wqUt3I3YsExwMH63IZLMkhcyfqdUrvmYxeYOpm3vOczpVhV/+
YGViKqAj3LH6cX2kNT+UCefLgoY/iHLhv7l6KrpHENexjlBAqWZQ/NbUU3va21tJnVbl96tZkXvP
MS3cLY+F3OPh4U4EkPbpLr+fme48QjOxPYFuPKLBestLGlGQ+ziPQcfNhC1zyqr7TIw6grfDlfXn
0snxc2QMXekRP2HZIPnLgL1Z41G1Wmwlm54FwMOSOLDel/OyOPrRc615pleQB3QAxFH323H3DYne
RqVLL98XP8/MUlSpfEhyvyT1xgIq88H7VPbPdj9ZdLJxzIplvOIp/l9c92+dENaCeXk2tPh3ttDg
Xp6xXt3kSMAYRKcVKEVwe8Msc0haLygmu3WTVxZ5tQYjZytWLeT8T4+kejcGZNJe3tV7g1XTgrof
RO1YiyYbv7ed34MLI4PHzUNlL67tANPNHC3uu5eF345Ow4BS0VUCZF4QBW8XCb9dW1geH5AOxiXq
G/J1q2yEAj1Swm9ct9BIL3lk9OaeXkB+NIYHS0b3I2ODjW7aIX1ui0+g8mTV2Cz47AmdpAzZd+tX
I8F1ry2tvBplNmhhrmMHj8obx/2G//8rZlVN6dMu4RTIY9otJyHPlt9+pBdoyCyzwvc29gE02u2H
w0MRE2zc9ilzeCvAIHBvIjhKO7lhIoohn1k98N7xAzlR++ZgbOKcOZW9elgrsL19e/ISjKrraxPl
KFgklPnfsXqGWRp7jP5ceeyAqUEy1ByOv6QgQrwGAXSonIAxuto/bzpAU8/8twDRcHKUXkhw+M9/
hzTtgUpuD5MBpKoH88fli8IcQ6YbrUckZ88g1U+xSmpCIgTvWM5g8KctrJ7OgcEyAVejQ0crJM/v
6fTCm0reVW0me7NEVqNe7ValMJTQJTBJ6N1ol3yL+R0ZjKLzJYE+ZUMeX80FVGhRGHviLnRlaA6s
sd+4D3+f+8E8F33AV8jxWxWxhHiPBoHSAbGfOPVOdXt8n+TMiDLABbD6cO7Yf8SrXAAwARkVlQiJ
PDJ7rUdgAO2s97QNhp9m88OG4bwwAag4O+tYW8TaabqfRyzKNiZ4ITHyWqQM+V2DZwApnNtPPHT0
ornViUlt/0mDcyA+V3ckRtQ5WOB1abdsxzqNNDkIMq4bne54VwaqEqO27Ru2lVd+WS66ws+feCbU
Fq8FPZQQgnJbfmaiuPAEMobxqAW4jndlAqPxF3+YOBLMJAZDC/xFT5JtXaAQ3e4YkKiPMIwzkXZM
Zx+IuJg9oIoqBnRHPuj7g77KCaGomMVmBbT9FreM4SUduiUK6wJf4HpNudLWyIncM7vBNsEZ00uB
ZlD3NINOHeEOmGLEZxxwZOpms+R5H3cqaLyqd9drjIlrosKan0FGY5gT8YG8ZLhk3DzHH8MwXgoy
En2N/ISiBF27KfohLbCsgE8t8GNz8Sehjmfy8fx64UgubdfjB0wQn5LXg040zNdFh2XYjLAqiWEy
MRx+arIHp1bnDnqbCvfVY+MawSf/geS+7xT3Ci/Dsrx8+0KizZAVaxNiMnEodKUI/R4rGz5dgena
yBclNb9QyVFoCEsIMY/5KOFz+SARxc4J24DEcXu58GAHddi0L+ZaJGVpx892Vqf9G/XZwozpk4Nd
dsfPuL+oA6uUWXhJ+SckaHEgcW2+r7sYAVsTRc5KGGeQyMjz5eBK0XA/PfujsscFkoyEdI5Phx+U
rPVEq7HtOh6Pi000SmBwSud/SCXXMmJR5TRE0desdHwp765BxR4MdxoFgDtZ79rMntTNEwGgYpri
W6dN+zmTpPTkQyG/nSCNBaD3NMaJ7DYT2HdQPuis499QsAdGe4egBQf5t6T3L8Hk2yrSOdG8yyA6
irqDI6O0BWbMuOxtVQHsFwE99rhC4yKRAMbJ0XdtHsYEW08cfbaTi3MBbpX4H571DJizvSQ70CPB
g3os7q6rcNqCeUOh6IzyZ0zvWzfibbixCB9RF/CgL9ptevQ9OxXQQ8/JiIAftizBtSJHZE1J/son
rqXmPPeWuwkTBsCRPjteXKC2Wp2P9DbmLgwo2l5lVAuHNZ25XkWvpz/ToBU0WI5nO5Fy6PD5nJW0
xRvZIq9FM5MNWOXT8/6+JJY7sog+X6RxEUySlNa6M4M+cgFql1QnKdsVvS3ntUS8ULxGVrAGqBjs
SI+Rar2ZvHQnypgeguc6IJZd5fmtlKQc79tJzReFOYl/Bt7F6lj+vTL5DUw1SA/lL2+1qLQIS6X1
6xaWP8WjZQBPjRxgysdWYTrLYNvM/FasScaWy6IbBUF1PalifZe9m79yb1O624vAc1j9H8BGhNVk
7vWUQjTealn1uvDVg/r4bxQUgFnizKymiFxe55ef+whLGrEWbK1gNUtXSQHwUiKIeIOgb76jk5kH
OuCzhcfKqLnhE4Yl68kH4BheF5X3HB5OHU33E6gIA3uhmjsMXCwBdnFIeOsa2SX0isEkTl5eXs1I
XzJ9qQkAEKO+8eKT34c83FWGceqW+C1iv+za0kqG/bq45BaPp2ypjNMJ/qllPNjE5/TptzArAhLj
W073qSpyvSVZ+CFS34pRy+isU3bbcsEUE6rzPOW05vEWb4HhTiTf6QpPk3s+HqdbHmCKO/jAHkPL
PQB3C73qwwDcuen7BA0YqXy22QFtWCf/8qX2ZhIYQaHvyl79BcyS+ZrtKFOMFTNQNgqvykrNMqEo
x9VVG6NuuuM1Iwx0tDuoY0xZD9JPZ30b8zaK7+End+JdeO5HacYlgmxOPZlLZdKHXxsv/PG7iiHt
/K9hD2izzuRs2Ik7Uo6V1aEKeJMoCBU0U/fJF549pjsK6mwkk+n8O5OV02RilQhQunrEpNq9ioFy
hq0yDpkJOBfW03QewHBjn0oopNqjmgdQJbRDOr5Xpc7O6UarTRx8vvuff7hH/+diNRlToa6vxNhb
MWsL9a8QWiCGVymoDh/bFEEopx9/c5U2+PgmVBsgEwki/Ie+woEppSbo6ELpxqx79VcaE5vTSXVl
U+QhRhS6zHp4ErDmFJFLho3haqxBas6dfKf/zwJ71q4ho+gHLky3ttX4pxQd3JDQM7gaRfUr60Rr
ZzqUFeQhqdFat3Drga+uORwciRwOBm/eTPvi10OvGVze73823+J9BtqO22ZAmmyqDQEtEUk4LVQG
IRSR5fDyDPBLap0AdrgaAqc48/v4Ods3Rf8KNVcIjGvcVjnm9dJEpHWJ9rR6raBukkVuPt26gsGV
YMpggsAeZCamTDlSHpnQpCoWgS4nUx07nA8VW5DOIQ4xh7C2RPz9r3mfnW7w5n/pl/qRwr/q0u8M
3I71rSnoX7OXtQ2mqkzlAaPt23yZFxCDeDmqsXMX3OzUX3OBLj8NYdYjA2bDsfivQLq06kku7sy4
tlx3x48xZPGc0RYgeU7oytbDX2DAIX/6R7V3dmN4CnclwsupmOJedWKm4ePwxlNiodJNujiv+j4G
kxoHKYdDJ1OEW3o1Ud5ua/Mm3k67TbdyHHtjVVqvqIZ4zqm6+uVTOY0mgRm2wa30C1/8wVmn8Okt
wxbdQVel9TL0myIVj0Ty0TDiQxfcwioeTU5bdNe6WJ6idSZvHhtyD3D5zbSssCHkx9CyxQUkUS1g
ltxBm9fnO4XwoL8QSHPBp8/LDhOBEOdI5wgJE393CSRXIdQNbRNUcel2IYIYGfDem883UPSgJevT
JZac2Fd5qcNvmBX+FcyfA4lOl8YZIzofS7jK6qSmQLgUOFd/s1N815FDeTlGMUEjJ0004qOK3b7+
KRghLTphOq3Ddcu+Let3PSvANNczdVq/CEJivuV56z3mAwCVBbomaS+Ucrn++N3QAo5LtdC8c7GJ
XaSR7O/9csC1Yx+npGAP7yCWwMsFxlW+1XN/zeCKXz03RYXVOZ3KVjpCCV46UoJCKqdIdmjFeYjK
PoPueJr5hB6GHjXZ5Tx8sBDnqUb8LglZENdilchRFo/Xdm+k/SDi5lekX8fCptcr23qPQ2CU5upT
/D38IpW5zjeFfi0quHPWgisjBp3pEd3PDhkJdGE9f3x9Jf0Dcj/kjWfMQmPFl7j6U/3NfhSl6S0p
ktD6JQZrpyssK0fNOaBlFxMNvewyHnXk78b5sOT5SCGGpjoj+X7Y84ijyk3pS9YTAYSnDLrL5azb
t4GnEJBxspv+aOBKb6YSQnePKyvRt3VqO2yMSL0bhQwJ19RX1lakKjnRrU/W7rw2Hw22mQX7gyAb
ZhUwJPMYhtiyl1N85WsdsSbGIZLn6oo1tW9i8pbukX9YnCcSQaFYUnuJrz/SMH/IuVnSPIaQm1fc
hvZ8Exgy+7oMyE6G3dpwHB8yLctc+d2n3YJ+T1Fyx3d9xpCracn3BpIFNYJCjNcuLTFPfWxeM4ET
oesdncj/vY9hMZtBaD5+2pQe/tNy0zers78PUxdafUWNQsz8LzDX2Mw6dDULMoQwTUdd08bRruE0
rc26sOtWkbdLuBQe5Apw1SdfpUs8k03w4Fde5gJemK1+WHH8Y3d4TmDb/HGyoQ48Eid1NOxsfn40
cYxBdVyLaLdFJXGYrFAf1C4seI0jbK0IXvwmVqUBIy3G04LKX+CmgVuP50ZJoSrTiXRpkdFFC2t/
BpTcm0WLIpwySLGbu0bRKwSnP1Vub6MDUiaI1zb55gIRVPRXjxK13nQySy6aqG1M+oUHfxn+c6ZS
R3TrBdt2017uIXzbvBn8FQZqqXydqjhu6yQSJNsRJ43ZTZwkmprmj0sG2Fow7tWy7J4/WPsbv8H/
hH9hj9hnOA7+0L+YdQ7UJLHaWJh2byZspUJg/UhT59SK/SXwo+s4cjZPE5hrC87C4S6+KjtYcUOJ
YR9RcVldScrF7VKcq5kFMRpb5l8FasPvx0Y8+Pem01EmzBP63X18nAZUerPZFYk8La6QLSG//OsD
l9yIYTPvpEcpVypjNE0tivkA37JfRW2UJNU/3xX286H3V1QEDqr4vG8ytT4K0mgoipElXtvTbfnD
fvUwjwq7l12Yby2uJIw/Tdu3on1VT4X6Nq8E8VNae6iv+jCmjECXKBQin6OnRntSFkAZ1gpNmyKt
bsO+NttoqgAI4cGnKggC5TwiVT9EmT97iqhD8x9PeuxesV7Fji+4OlowO+mNNHhcwN+UO7baJ4Um
v5V9vadc36St2270X42nh2LD5a+dJjo5oESGABktbiFH2d96ejNrDXGZEhnbTJ1A6F3rPD8dSN0L
b8YjOlKTagsDMrpx6e2O/fELUn0DJirZKCffQeaJ6lbLhhPh4ENUZsDnqDL0h0Q7Yco7FbZdTbMb
NCbTHNIl3nJKIS15wnLrUEcyvQlBIIndoZqnRpWfqsWuAnldacqwq36rWB//doWltuC+pdREggKB
00BPbh9lrFOEzXAY8B8mMLpTxPBhdjmttu1RGlkV6C1xeSI90t2L4CyKtFSD7K6EN7vGKrLyvffH
zLJP+8JLHFDA876wj2CDuHiiCkEGyi3rs0rCGjm4Plmd5CktNmY6g1PmtfUK44Dih3B8jMt8QROS
K1hicRynbYlzcWj6nFjPTtK1ZuqbBf1DN8A5ddbn6GeQ/XiOH6mD9nOMQ5FfWdES3cVF+onc5iEV
Pz8ytsZoNtrkRGZ60zupZ8NVs2sSZKteDM2CPe4cC/cGWA3O6uDM3MtW2lAIbywFGE4i82kf+pdA
BOmgIIN+TKkw3bm2dVVi8lZj+Lx+LyAv/6FwEr0Ei0Ob7HhCucqhQsDuhSoCegiRQAS+5Tyozdk1
XgHjaQ/NwjOM5crYYkNU+dmNmuco0XqIJzdv+D2GnSJFfAxLZP3K9iOJP74oJXZFehfnbLfaFega
NYBgXe7eCfyI6roySKcF6J6sS1JgfncBpipVgezEFnzVI5L+2+y8zeQKNLtWuzET2LPJxb/j4ZCx
0K1N+3tPBBJWA0Ia5RRG4uO/TqW/CZbLdIZYd7P4n4zNgrygw3Uik0/NPorSbRsDss3P9Em2Jd45
5NNq+G9hKPJJFXHSzSWkI24erkohTqLZOHNfrIdc8nkiv0aTFI6ZsJmpadlQUdz2YyLJKOMJD0Lp
nzskBdSvcD6EtQaL2DXQ7ErLu6bAWbHStfqEgDd1/2hIft/hOVd+A58BHkmVw9C9vVqlAJ7IZ2Rp
GvcjGnJEVQvrKZhFf1rLKvpb4oNgUc5NtENZDmRcINaycsqJ4V4TU0YemPrMRrTVhQGzLLKS00TJ
ZjrbdOUoPRqAzhJgygB96FU2UiJO0t5eroAXA9e/SNuHV60K64bb772qHsTh2fgPfIkwsprp+mIC
g1ngneCdMrgtkq/6taMqUbdV+0uUO+UwX9FSBHpxmZVkCFg+l7juGgbh0WGjmB3SFvirtGUbVTXl
xXBFY9GtPWOMvGfEO33VXzgQ6nqhYJSMWomIel4xWRGkGVyNcj4aseZzaGU7BJpHhrfkTeiEDWYY
MSGfoGYTras243Dg+7Fhejv8vVvvaDQEsHFiDk0gI/Ev1diiZtjriZmt1uoYCGgEl6GviJQV6Xko
K/Fn3QLXu/Wp7lw2+tm53cRyK4DnIe26LC5yrprYoHoZhX4o/hb657Onc5elYcMIR7B52wJmMJeU
iCKQ4xgpf0rE+EIEQKlI5HDqoj4dnbq3ecK+2gd6n0l6czjE/RzD0+Dlys/y6FPVCP4tbuq19YpC
jspsEQFTuLaTUnAtiaOPIaTtMati8rBqqVeSjIRFd64bA6gNjehir/A7nFk9UoNhCDVWjMKa8xO0
qUENcLDQGWIcwCpWgJhB9kxTnYmoISmtKKJNlAupM2tUOUn2bpV1f3GV4CcSMdbS+sk85tLJBbof
i6mgZiGhwwVf1yug5pq0Koc5vq4Tyfi0hQNacjE/CjcG8My4r34neiDL/Q7BDBlzRXcFLjmZnX3z
eSlHY+kwUabq3LITUvA3jXli/RvS6PGzB+mW5Q/uaRjbbm5FexDO7ioD9YQ94X8m8eBmVFd85Vvg
XiH4M/CrgiDo6iEo8bIQdTqeD5EMy7DCJK19O0MKTsSwwgNBcWfd68n9MFwsL6hbno+60BSITIyz
564HBgLcd6utVVDOV0LpvaUuwKZvMpvNMqBi/WZmVaz21nlcQHBSEcTMfBvp0MVHyfBX+5mlheBk
DVEk6TLfRnG6vpuqm5uiQ7gDyv2eFyEHk0h+fm2EOk676KeX+KuN9q9uphqop99YSsZ2v3g2feAq
iQ5L4LWONfgsdBY0Fs0FLCdel+XjQgqRvgDOVDmfeOZ3eh7fJvNgUyzTXI9DajXgop1ohNe8DNJo
sjDywrQrR8RU0FhRjxdybvDA5hBAT2DvoFAwgcaZqzFaxBhG3Vw8QDQvI57XfNEdtN1DI9ie1j6C
D3KUtRH7CU7B0UP5BEIoM0XLfv4lWXrtWQaAR/BIAxtxi72AyIpmm1PLnYVGikn34TNwKgkHiJf2
i1Wsm0FMx7Ak1WL9Tjd1ukDAb9Uu/WLxONoSTmVb0gyoeaZA0KN0MvVXiFoY0ihnqF10dwwgjapD
gSPE+/0+DHhBqP8p9tFavcp5ceaJpZPJrOna5l7mUy/z8Yg22i3oACxDEqM3TfZFgg+5t33z79SZ
Lf4VYOVgMDFhlwQxAe7tZX5cHehEXVsIwppo3DhEunm2QEKpK2QPbMX3DebVGoAh7gx4RxJKvuc3
D3h5hC06lcoJVMFzE62R6PtoNIYwaAUprGZYsMzNghx3n9xGe2aH0EAcy0767N723AnotHoMAfpX
4uw6XtLRpRJnICKO2wDeGqpvrfoDwbuV/ynTT7TjhLZP2I62I/O7a64J/IkViX+cn2LNUn9MPOZr
LCSdgURa5KtFDlZ7+cA3wAKmvr6Rp0NYq9FUFo3vG4M2dnGrHqQn9MNfwB4B2UfyOwiuREooltpP
SDhR5wc1JKqoJ5V+0fPb9qOaABhe4CM6pIIbEcuMK/3weXQGJ59zeoc4jBo3wmlMHJ54H4rZ1flQ
O/SHcS1HUwFtPSKdY7kiXqFlSYmLdGYnoHBMwIraUAFUKGzUC8WXifStQXgt4BfAPsMCIvlr8eyo
8nZWVtZZHyVXEIV1x1Y89CKIODBL7NQif8O/kzms83FkQJiS0SMMGBPVUEykmj5NPw2Y1axWo0Lx
fe0e1qR0WBplW4Gkl2P7oni3953aFqABRHggAMRr9jwQMAceFkpU2sNk7GHgUhDkDS2StptgQTIG
i3+zUaezGQCyQ1keWnxG4i5x5mN2u6ds3Ud25sZZ25qIrwBAzb8A7P1xlM5fgi+griDayLK4pwC1
guirAZuDXKY5IwAzzRsQoUUcTmZXJy7h780HXjEg4Uo3VD4w8SjHXw/BBSBCixoBUrBoupBb8USe
E/cOekl2J3pw1ViFLgG28amK1keEYnBxz4RHLTOMOPhb/yxDVFOEqy3fcp6zmBLWLso28XInakkH
nRNHtTjnFi2znybocDEzBoWKpMqC676wMuAz+J5Ecnjpwx80vXaJt5fhq5VwSJ9GKXS0mx8NW+R0
jk577ynYNHQctA2sS2rGoWl9wbA8Vc9oS/e44ZUzBHOz2G7TnLRxZyDS8YF5+3f3piMW9DFudLbP
DywRrjy1zWhq9w3NDnRjcYEsDeYwIscRzDVcG87aW4PXLphYiaV3hrKEO48RZizHfl81KaN4sopv
W9BUeK182BA2U5soap+F+N0GZX/cySLN5aoCBBki9wIBOGuRroKQEwkeF7PC9gC3mfisK2/KBP9r
2Knqp2g5s7+ZynWOv9kzQudWpI5WKESjDFWgBO4qz4+ciIEU0dQSrKN7x9s5ULn6eH7wIsik/jI2
/Wvh+NZjd841ZXCm+OWQGbHeS4s34zLmzNnU+WsBKRgtRrgPBWSDnndo7Zdik4lgNrToFCqdIC9M
L/cOzKvnQjgChcoBTGObTyj6RiZxkCmkNJiztdq0dcsebn8jOwX75nFZXTZO3QmKRmdxMuE1Md1X
ynWeqSOhzA6tI3MAZ5Q2AB3aO9TduMUVA2VhtU2DOJmnVdnQ0zhsgKbBWu+9iYsT99Iq5IKppRN4
ghLY1fBw8cPK5xjIZFHhUE4bK5/kj59EU3w7tmoZw+7txux1SpwsPMP1OI9tU0uVPRuSlv4N/8+V
m0dHcK6GqhYAa6OTs+SfvbS50yOHbTlx9GNZ8jybSWTikEGVkNuTL0Y2cIZyrqxZz0JqJSgmV3Tc
7OXvOUuD89jhiv9UqD07K1Y6SuSt82XjdEPp1PRd76EZx7/NvtY7DiKgrvqoe78n0b1B0qNJelSU
1nswLcPkTdAichImHF+3MhYzUOt6OSMkLCtAhy5fYeF1ENVtvgWJJs25zgUWj8lr7lc/0eEvLZ2I
aIfHVzVCfqdJvq8qdmekLpSS+oBQ3xKXAlnDzCC7M+VVcy+1AoBaIpJxD60Jp1e2fEPkgq6gYhtn
vufmpHQrwwVw2focPfveewIXi0JEnHVjf3BZbi3t2FCDubK4gqoTMpeQOYq0fpEn2Ug8dPFsEGrE
EGQQ4HN/D4QQ4vIfLD+WXD5Ocd0abh2NSXj7VeLxrs2UIfiabbu1tv7rhfSZo9TumerGxGYdl01v
mQ5cQ7IgYGSS8u1W/kw8Tkf2mq+70Yt4XtoYkNdk5wDWATswBkK17o9iApYumbUwYU9LrvXLFc7T
VUw889PkQa9PzNd6o6xSuM9fc/Ve9ct9Z2uhonnnDjv27aGBgzPaLmA30PL3oL+/6CJSp51DlZzo
Y/wnB8wtCrB5b8YzQDbed4xSVAvRoAplBidKukOBZxBK4Cya9/KnXWWlLESu45sQw0yFyng7mZ5g
6m7j03zUOLpYwa+vgoK9YIsUsdm5Tn17fyr+VL45AdUGFRhKw4Ot16X5Z3MKjW2J2kT7OwFaNOSg
SYfnhOXN2knevL8THzEoket1lWX0tMHoxJQHXXJevbBZvCd4EyuFdciX0RHmnJQ9dJMzbugSrKEC
TGZSzPSndLvvCt8SwFpLqeJWlArYqKFDjgam2ks5I8lm4gTZ4Ntod01JewHDrEFH83zuyXkZXt06
rfAqpe2uwr03+MCZW8X7mP2WqT65wV/msWhhTomCoojBPvPT+En2nlhV3ZWyOne4dPFUZQnLWObk
ed/mxhRL0Lt+//qiWW2C+QL5j3fq1VfCd3qOLQsjm7MmWYMvWboqvsL4xvUvlWj51nmm/ChQA3jF
JgaTDT2EmVIzNzbu6Pad6sPb5VHPMx0ndKa1b1jHnuQSVUjbTwvrbqqCMD2b5tUR2YSf8V7yTGTB
SgpQfbyTV6Vi80XZwCFcMR1fYneIX5JsCvWAnC9B6ulr26piV1KcewdJIxQpRPqqIyuUvBqlAb42
HwgViHoMzAEpQt2q97/rioxxe+u8OiHevduSwQczBnSOWUXia7evGp0/fg6I/N+YIryNcf8qNbpJ
Zim2O19ottZSSxtA76dXGc3+727WAkwhIINb+KiK3hKqqto72LebILHvpwkA5i0/9I8iN2Pa/5CH
HGBf5NEtX4vDRDwmiNiCNTrvAczPt653XdYARaciLZqxQBTkDFeBhB5qbzIgntcOONO8jd8IgPyh
65NonyMhjwYLBdNq6Yjg3bKrqYj821IuPYvv5AnUTui8r3I6kOPqsrKRFg3ZOmNlMZ8UuHCoUi3P
6xZ8VrzuOm4C4GaS/slhWl3u5LO5BcfteEIk5GXFx42z6jmDx1xlvTgp4qkCIVk1zhUVKlMYDFYj
BqbX0OwdnllUGbUehTwjnWzlMxkBHzSD4le2pTsYpzSeXS6hYyPz7BGggkCkqNlohUNoX/79hFZR
pByE29LwPOe2azusVBFlOd0R/Vx2fvDwHGmgYNGBa/XV/RuYzgh1aBRAin9cDUbI4sKxqVlJMl64
DNPirJaTh5WeKCw/FypytJT7ykCVmZsWEtZVQCTWv8b8Gy88EM/1x1IUwrdD2WVJtkNm8sx17bAf
5UDqph79THdBs2k3Fi+XrD1Hc1lUczQ4RCXvjcorZxhQ1+ikyEK+MLuejOEOmZ4dDwoL3/ol8O21
JhC+LdNu/YuqsqN+GxA+1dtguhJd9CuDd3C6rHK9ahMoNl5aesPZUJh/JZUY5qI4oxUCe0ahp3yj
LPYBK9N1ZmqN7R9holpTyM4Ds5Q/t3EEZKakik/6p5mwm/W5xVZZy0JRvHJg9Df+u30sbcg9T09K
cGvwJgiyz7EiUc2ZnQ1jqSnWzo/KgyBAYDrIBsAazjxvg0uBKteh3dc74FhMVAP5UKaHSw8unPz+
DbL+aRPW/4fEmBLtUCf8YypClEpo5Ymw7zqNzDwNclWhbvQke8DrjdW+SoeZFOgQPJV78Pmp6Ry7
ACy+tc60VdfyLYONfQM8VODT+WzKzay3N/XrNz0b8boyBoycm6HgUK5DLhLj7pVoOwBltdiybKt1
hiMh4/3L+YXMNunIUgNT7Oho59/pDId8JsyxmX5TR4uzgoeZquqldM6to88Ipp4oo3ixywnSZMqD
CqXD9mU8pPn7VYEzU2PbVC2b4nyMibKpl4Au9n+8ckZDyB5zlLcahgbyggDXzf9D011nAvWjgEo0
eaU/g5bx3QqDqkKtPm76JkOU+Fg53ad7smNfqoj08dfRLg1QYi6ZoNeHcwqLakDhLzMKZyG6rGFn
Xd68vJjW/XbYbSFPn5zUvpj+hY/4YV7LCuwNBUkAOni+fWOV2Y8OWlxjYIud2HPEOWUdL3fXTd3o
bN1LjcYtKQuSgPo29Tb9PtXXgji9A+pNLCNjtOgPIOWzzRS1tofzFANw0aiP8pJfqeUukrNOGmKz
TUwDH/LnFqA6P57JIK0ir3KHy+CKm2tU68CxXKiClWcwtwlFO+z9TW1drdh/sW7xspDcDBx9awo6
0YMhpD50ZcyZhg7hOqKw4eeeibxFxNcQEn0bFzEzMAp9EK3b4wylzjPdBBftqDOQYBhCPjt3XXQH
ttu9/vtgHtDMkMhrc2tZ84DnnCE+lYdjlOMtgsOklkm7dD15KNGskQgBBSC3qCsjuS64WCr7K8PK
rqXeRA4NoOElUQArsTXjoYLaIuq+dF6GzFUG/ZsIvHtfSdYS3eDpCRSI+ZyE5GcK97AxcNGJ3Vvm
t+lCqKgKE+anSc4f86ocmTu3Aln8M86OGu1zhS9/2MB3i957HVS2F7nBhy7zCx+cZO49Ws/1xHKC
SUk3/dD2NNp4RJl/SonI1jzDAwI2m250XsZgNl863kJR3uCIoYyxy2gDCV3HPhOV6Y5khRZGaMNz
bjvKUbFCn01ppT/Z4cnM4IR2a6fYMybG3zpB4Ny63Td+LMEgYY6hBUs3LZYItMTH0C8f85jP9eI6
1PSwRGmZxLszsGRTNl8evlXlK8JhpBfMhiGPu5135lqjX1TfeVEFVAwuwUmLp5+z0OoHWXzjaNiT
ZB84noSIoIgcUlk/9PG22rRqGMDwZT+FR/b2zimrVp5bKtphPtGXzENG6UhyKZcwpEaaOG7Hxr6u
ypX9glQJtbHVB+nmjMKaGhInSmkDiX6EoQIrHxo2ZzCcjHg1pN6WtxmdVfXfV5IZGKsz+BDBr0hP
Ki0rURDXNV6LOyD+gY3hOUtsppNoH95u9WVUgvGkFs25Eyw+KufhWVARBADXLWSyd5LYKz76p12A
DIjxtkK11AVbrLkBvi4rmezrzskMmAyMFosTh3c4No7ZavXieoTBif0Q2abaQPaZHZi/fVXmZbto
gWJRZ3x1U439+922Jjk/XZnwYB1xS41QpLh1ZzNUS4ZlYlc64tQExQIqNgZ4ZPWv3pk1QjswDIaL
QvSxNeLlEZTfg9E1nvRSD6jENYmrWT9yWJSjD8WTPbXLjkWAzbkT5wbQI6h76a3I4N2tZoySccmo
2nnjrmUcIzvAX+RcoaiRpA/3Xa/0nTjJsjG4aXSlzpbm/mfIm09Jma242xVzHiX7nMnh4sPnjPkh
+phBGQiAlQ3qg+WnzUT8ouwIxZRt/nTo2T/Fwm/jjYNCj8z6bxauiUvo7/d7HS5hLvimZvvlAv//
VZmm6oFUDu24uYYCvm5wh0YUkluLIxCup9DdnbdkQvE2LEp007O1XmD3ASdkK8jVYSNAt0pNkyfy
9g+LHfcKhoNZZ4TnkBY1+LC1yPIyyQg2xlPeXmMGu62OYhC899bv162CGqRvFOpPuocpLLq2nKwH
orn2kB/JjtYy0TJCIG3MZl77Xsk22Kd2793OckVxv26chMkaG+Q53wYusNR3oNT13tXrwmt7+rd5
jPRHbEwmDHp9Qdk0SPcib8G4SVLAcRMDMDnksL4mpfzdZpvx0VkWHoWG6zcfB1ryneCYjA0BPODq
1/ECC7mvy69HHcSBWr93JFwd0xBvLkIq8kqdHDOe5XtsaCSDMBV2qXjWugX8zKi2otNAgD6DO9D+
SJIW1/zGtib/Trn/AN59ftrlP6W84uIiD9w2t/Uhap1dXgtJj2TwNjghbsopA2RbPvMQuyswPM1D
lcUiM3oCIcmY80YFA5vmctMnBkETe+x4IGPUQ7pmDDUHkKB0fTjF8wxe9BhnMiFC6k3yamlXcKqK
DMNBMMamX/DBO6YxSJP4gWaEHdw55EtpKUk+x8iw0DzpeVJkRA3x0X+3S6KStBInN7d/jSJSOIHc
bNIlLuiEvs+si20q7W72pqWDxzSiqMRHvSRZB0yDvWURYmSfLqvCzTMWIcTFoW5ay29uASWx38Tt
BbZEyXhbWaV7p27Ju58rynHQs4FNk+EciV0EZVI+VLFRyRCv9+STeTRsQA3BWakRQomn0I281tGD
HdD0mkyvBATirjnjk5qUTjgBZzX7rFUPrHQIygKm5fDpAT9FYceZ6fA5UD9LHHcyOct+uMQFDEy3
C3kQrzNlTEj0Q/f21ZxQYaJM8Uq9NjR+PNbUHECl+eDoFJauzUGMlDZicT3fiEyidSsuvLEZ4jCv
sgvMJtyIm36TdX6K+FFAqmnh70g0xNtBp9N6qHd3G/wIBLoWZC63yTRJYRfHeKsKurig2fpXoU7G
8nebvD9PwH9ZxQeLtMSZJSMpu2nDgq4zyBLfk3eaY3LXqdI4Wm7kbh36mUosu7EyWQDjvaUHmnAW
HYtQSD7nEPlw4zkygyhKuzIChbtA0gPwk4/mkKIyR9zsMDKEXlNP6oVzQ5AdGpSvx3mX3ZlXFWAt
NG6TmoaNsnbQ3FuPQ2uUT8IyDFg6n/FQ6l0OA3zuyWEs6+XBRMrVS+x1dzmddzOZnfviBZTuFsrL
5S3RHerSjZwiaGgtrtoF1hdxcvnw1HV0PmVs6C+L2hzZA2OnwQLkoZOcHR+Bj3uxPHSnKB0AF0sl
iftGV2ATmL1ChUx/WNpynyRdf8tbhotx2WfEOSUPXYg6IPSy5/fiAO0yyWDK6OIwK5TlOLzKIM6x
Uh99Mm8pdWl/faLpZsRYrIPuwk4wjkcU0W3XBNpSTiDzPjlFdSTFJUIR3zLS9a86LOzQ5GVHjLi6
97QDfA+XNcgNzrLVfsnAWSo9fyNe1d5CXl27O9yM3GvylPJ4fHwEHhkzqnZBGXn4CZevdpBbOs/Z
f8vlgjwi88RV5nqDmdn5Q83RA7TCDHMRJpjFVKImvj+4wlYCyJSvm0GdrUHWp05T1c76u6Rx9hYQ
N8sYho7R1fCbQ2m4Clx9NP1cwUnQ8lRq60G3rTk3ZMmfqLv0ck4FAPCtyNzVetWKkvPh0DEipRRz
QTz/6Nn7eKf0Hirvro2REmM8Wh0AlkbgTgjzP9wnn2gZVqRh1QGsRFCSBvMEZLcbplIi+jojTOF7
onE8hc/xKLIcr0UyV/xM8nSCRnZHaaEPxJF5fY+Mege/JZ2keWxfTjAG5O6OKkG2Zzo2YEQlfnae
S+l0wRZUPr2HKvWs2hgwKXE0Pj8espynsKTsurw7/yAbknMLuh0RKFub5HXJY6mmwcic/cFtPbDi
L7Go0GVv3fe2r4sHW/sFnnCwc2JgIjaHYdgr6agXMqk3SPpdzImC6L2R8j7/Q94+1mo2oQR/SKem
bPG/dqGAyymV/P7Ib/JnVTgCv13yloKqgikHzGsOXPoBdEuZMfDF9gvrchKp0JnugHRkmPYiY3Bq
DtxyDTgl8eAP6yT1mpU5ayi1SQcLzH6R9tUw9Maw6Heo12nq5v83TlTLVagawdkw8qtZnqBghYcj
wvgTkzxdgAhldMydz2P6AUlSslmF9bR0DvH9slMKd9CbfJfVngAgBUQKBrLPndLH73ktfHYly0Cy
rGRV0PjIPPUuir0ikFCHUDdNkW4QZNELZtb87Uf2UmhmS0qAgXFjTrnEBRaQBqviM6r8//ptNPn6
VdtT7BSGgLRSkS5sRxKJHL19K3DZQ53dH9UgtydtLLoU7jldTHMxZOZdlCGQzsGSiyesc1w0peg7
bAKYgY1uEsK1xn+mz9McPPZQdFRaOp/9QJMyO2LfeQoBxjN6sb/m9r0xV5/hsbxY99ewtR31sMrE
jcYXqkzIVvmlCehjdVPkp4MhuX0ianixBzz/1q6rMlZ/4ghqro1RbzzOJBw80LZV4eqZ7wpL6Bh2
AwJAA2DMntO+T+KFv4UbjJfGH7W2l0ZuMogcvE68wEGezTaun5nhBs178dZpt0xUqTnPKFV+58TH
2THssMRD/m1Anv/Z0YBH/hYdWL2mkV8nSfafSUBIqZ1Q/qwkBAd805YiIoIPUuGvxeif4oPsVQky
cNXYix+msJtUAlE6CgnY6sivVTK08dKqis1eGCzIPivkp6MRKIGwK7khU9y90ijiFBxaZGdEzsun
a34ZMbLS1rzv8J66hurxG1fdUaSlLPXSlfAmhis1k+Q+oElV156P2Iz+DARuffIsVENQevUXPk2h
ReGPrkd6/fHhawQX0YMoOyRj8pQokRAAIISKIT9xD6cvWjkRiWvAOW0jmrdEfeer3VY5slHa4ss/
iAGoHNSSvUbRQBBoTISvdkFr9/4H2PzZTNOojYUqJXkIeKuKnrxgxKZcSs5kIBravGe7qdS49tFQ
jI6MjpEIZeCAEM+bU+1/Lv0qEj2DJHMlDMJL0s1SUY1sir8LPdEF8D+Uu4sjuV7b4SnTacsdwhRH
CxAEmWcFqQABvBDNHplZj2Mcw9Ryuw5E/6DNTdqBw1wTZWV35hmYPoKfcdSiwtPRHK78Kjy9cbxA
x3OXI+EZdUtCDKRbAgW3Qey3phONGJeQ8CR4N+kXS3oLAPJWSqkEQclK/36dYdMFoxKBURC05Q0d
FSAjmVYEWJmB9J87fByUchZL2ru5bkmDIllWxigCWpx1BhELInAdXVkkkpUryfauF0sVwvmMtS/k
amjGzCWu0P8mVSE3pdDpIH18zM47xNSBAFBCPQ2jwebwiAQqxZcdqw5dnPMZuglbdmZDk5wrI6Ae
N0nUxYjs4ZqBFdwj6yQu0nKFypt10QgIsT2Obr9yrN1WEVCwlMx4wBFwsANOTUOsP1B+6RG+WquS
9RmWLMp5fhg93hfEHwj237lOGXzwIjEx33cdbCvHSd2b7rbNhsA51yVWPrupm2tA0LLQf26TK9eu
G/QoZofVvpi6NKF0+Z2llOw9eJqzYsX+yDHYGp8RV1hEunHXcoGb9rTvt1j/0j5uen2xV+IU0Yz3
1A1aVc6+hBtyqn3PUXLaduoq7g//JMTCY8qd36BphwQoeziJ9ALrWB7QrRA1f5jmvA+FH7Rt7URI
f7WlxuveqbCEz95VBrWN4ngluB30XY2NvGg/fYhEQjx1E7AkwJF1ORwnUQnx6RCJdkscZK6aPKdQ
JhHqF1jR/5SuWm7UD5DPVJqNzj03sHWDbdNjhwR6jQ60nPbqQX/Y/EkP7DarQ3bs2honG7IW2ntB
iODsNkM2IXUOufyzmS9lUMftrPuj9DgH+I8GJj7an7HTvutFaEiTHxExfJmAz6u2KRDhRDCpEK1B
JTGj4R57L7NKd3MomBsXPsgyCijDP8Ky/+edcB/MBVibcKnLxoZwlmL9iSdnXAle7NarXf89mej7
aKM3AN5P5epWPrUEZGj4AX+H46pqGWFBQJBBoeuPBgjCw/BCmv6EuRmOlLi2c8P6sXAtTVTU8hWQ
yWYCqj+rB+3cuVPdpbgOnvPRO4pzGgqPYk0SV8Ca5SCHL4i6VvnsXw+TC06aiznrcv3ezlI+iTZc
JzqiUic4zaHsWEtsHqfgPCUHLBa736DU0tAwOlAXJSqLZQ4jgzbPmZPzPCcPbJ4D0P8W2nBNbQw0
GbeOYIMCz3bbsWCIJEAAkeD4ysCMTRF08d3XMo5eHU513oeoYR7iv93oiPG5J3ma5ISx5g2k+eEn
5QxZdIMU6/ACu0eBRBvGgTS06MALkZMc8QOgEr7L/dpKeTyqvj6zo1v2yVB6t9Mst+NRbmqqUNb4
ChOvt/o40wkFW48DqxysX955EIZEyXL25qFnPSctLu/5kRyF1cx6Bosm1xk5zitZgDRQoPXcMq4p
coK7goB2VcCMoQhGBRnGM71JgfAm3rityfQZSqZzhhbueNSkLqG5/nxsQDP8Eza9PQ/GkOEq1QT9
/hWZJEXikKUUCaAfFKOJzQHDv9D7KuPgBTmV44DnUWRcsIfDjxHJmUvlEqj8bSruxErtRLgZR/HP
VknYLVWXImXfxXMs2PrLPSfQ/xkz/E1iUfiIkBM8djpYQhp9HovJklA4b5F8MMOFx+U+KWIHZn7u
SVPzURGvzKZk4rQ/cE4Rw24MWQZSOvm87k3TG9nZyI9n0APla0tCl2iWXgLTZGsfVtOz9OFd9DvQ
RxEr5CAmLEwstnh+m4Ts9HE+DpX8Butnjor2C6hTrbgsrVwjZTyLlde0UCuxibJ9T3UcGfshn2c0
DvbLOq9fP+8ANJZGOGq2mQedI62UisW31RIO7XD6H5cgmwE4MfMCX3Io5MUTXhUV6GWCjo3kHtKd
xnXa6U1mELbjB96df2mv0FQlmZ4S5LrggIWZEIDY+f9yLIc7MHyQTrkTLwO5h/cWgpUs7CyE+NJW
TzSsAooXet+D3Khu8kfxcGtP2cI15mFc1MLl4TR7gHtoHQT041jKF1VMXqnIY8qxCTxVy32gnDtW
aRUY01+JmDOBN2hvH5WlqxR28GvatliubuKobQ/9EAqSA0zPLUWu69vjB0fpUqLQ/MgseotovHRD
hKEp1DXuYu5OzC/T2wpkG6IBuwIki2Y/yOcWTnHseXr+aycON2/dv99JWINxTDWLvmT0Dg2Hhfbp
qaZ69pio8f5hjGtM8LOdH8Ys1cJNQ4z5FPYv5mK0+fQfkzdxyMC76nLCCr/ah6vPzeCrIXvpfMPq
ny+641ODlaM7AdH/Rb1WKnTu+wMhx+ryaDosQOTBlPlgTJoQgqx297+JOX0cRW00tdIGAVx53gtX
6Tge+uKgggvscgVZgmIk/D9/Jea1XWpaFEphrHT/0xsVvJEFK5o/Ej+nJTzOPy4Uzo/HJJDWeWju
W2gOPZAeYj2yVDKOZdS3lNgTW12VNXbqdJgM24nxXHDSgQNymoL27zDIu4Rkabj+dbcYGFrdHRwX
8r1lPZbe8SgYW1bBHQk7A+tVTPK4aKWBe6FaQlr+VeybeRoqfOaynPmDelQC5rsNSqrQeDaxTUcd
uxRXlwi+OPTAwUupdipsyJcnbhLsEeYCdhEnOjSjhHu1eMwp2i7kMuq/br1anPeyiAC8j51dxT0m
SgHh/XMPUrD8CM9VAZ17phsAPl6TI8fWHAKUyoBzG4pyHZoA/jJuZEAA/j7SKBWWNj8eXjyG4iOM
uJ8iIT9RxAxN1DpO1ScbHf9eWQph2q2KdF+xknnOTw8i/KsnMjfyET8SHqURJ7KPeDbzYaMlKnkz
djhsh5KtJz4jXEFsaMCks4l7+yKNAf7XgLy+tTjoTzLTptnoq2CXeVIEA0J1bQkDRqIEmjmH5Qax
PItZkN4xQ8tfteq69vetiyESK5QuETA8XDd083vpjV0vj8immFfHadIuPTGQyz7a0gMKgJz2usAN
bn39/BhwaOebezVtuI6yP2cCLbSoWoDoZUdmCZmQOr7lkq+j5mP4VwNNR/9wM5Sm/IcRTPVJD7+W
aM+u+R9sEJ/Orx/T4S0iXHwtFpUQ+d3cVAxYrRN6M0be0SsA9tbG3To/d+eeyxy5w29kxwnoXq00
m5uIjbzs+/34ATebzv6Lsn3DU9X7IQraiyItULoOjHg1xtyFO+k0F3O3Ue7PauNa0CumDU1s+SCy
pgh0L5uDLDF+hC/5W+lCRZwOecHxZZgSprqIgUbpcceJv7eoU2os9En0ABPA1QnIfcFeIVs4n+Ot
u+/WP/wfEe+1sGMbrDeQU4q75LXQVrg3zSzvalAANuFUG8AjS0LxpR+HICaD/GIsoBkVCnwQtGbz
0PABZadJxJqBhwvWU1klcSyT6v9qX6irkq8XCWWmjvsCEt4D6PLrcuW/8djaT+jlKBWwZ3/mjIB0
7UZMSMiNo9WWp99sFVIH0haQ+fk9U7RY9ylVmTaRdJz7zUXhCviyTVPcGkDY7j+WB14j+oRowfpV
92PQTLsjA/SCKka9WLUrd14RpgdZFb8BcZmO0UQotm+B38pS6jCZlWdxuGsqHSbPiy/dUEmsposC
bI2RzM00jPlkF7kmGX2Z7J2I9y83ZLEzkGOcqiIdN9cL/Lw/Wc/Y+X8t34UhrqZwe+P2uFJcgYDD
HxzVXs7il387A3xc3KBK430zxD8ljPVcCqBPE8Do7kB/0aVmCUq8SUcrAS3fjmoXMP4Hsdoo54E7
EeCAIe4qHuqOmM8EOb4SsVvv202G+PEZ0ZAdlS4J/fVXp5/FHF1f9RwHG77dGuR0M3uhxEu3y/Do
t4e6Dix5xaLKFcMbA2Ef/dsots0L7T4hfJziKRYC8rKYV/WbElP+oKi1Tli5RFgHWBBHwXMa6ber
Rg2NgnNb5hEXXtxwXIqjYkj+Jqyl62v+SoGShdEZ6kmrhanxJ9lxu1koKeQPIU6Rb3xHANQXUtHq
C5wWXcznIhsoc94voJwQjQkooDqGmXX9xlGPtXo5o3UzZtqTZqd4Fl8itVlbssHIEJF5tZaUAcgS
wvE/4mrnDAh+8ZKJFiNakI21jwirWKh/9hFroPM//EkUdHqMOxWSoG9XEQc1dXVn7cTIcMd/E3qb
ytuIp8DaP9nmsd8wExTgU61wtIfxfr0yHmOBgqamS62xjHjXt6nb7Eva/Mihv1814wHFABNbXo+2
Ax+BMxvyxbp2ZAVIVrBdgZMZn/Ncey8Na330SoXPnn1XL2AfEMu5/j0JmNdqjlq9lgFZ1amVwNlD
Jtto96KgsLgOcuIQtecn5ydH4ceGx7dBpN5PVKpDA2M00Lobyr/gk399vg+QhE1ou/HHVG3KrRrn
28sd7FzMlyPrA9MwpHa01h4unb+IEOaEbDwnqpP8F9F/OD4Mwn9FboV5Snx9z5l88p1wULvcRUOE
7TjoHu3m+xMclCIIrS1rkvotvKYH9uv/fzwJ9Q7eyKFs2Zo4P6qYaECtY+w2xHY1XmD3vIMVQrnK
SQL7+j23fv/JascqhSzMNoxXAPnO5Z9JgnIJr/BbwGaNXCz3Xkevrnc/YqfgGsg13pIHtaHZsfxP
2qrGGrHzIC5C4sIQy86MOVFbyZzgVSYOQmWLp5m7IorQ/vdBpfghiMaJ61mjPtQ8J5H6z9Ur1rAQ
+bVWnNUKN2ySwy/OzfWy4vnXUBLDg+QaVnyHlckJ5pgJW95f0chauO+r0sjzTO9SkOJc9BA5vCDn
7f0laKLyDD5XMQDs4dftd9MQ5QJA8vYsTEgGVGoynGpiZeWLziO7TGbKwHRql9NNlnH2jX6Ufq54
cyXTkV0x0FVghd+6hd+cC16oqveuMrLTY9jaJcNZkkrkycsenXBa5w9Bb3hkTRmqZnFAd+T4aOD8
kYi9FzdZ3k8NPeXXFAgtrVdC5mhaI/BC1masQobUAN9S9QIaPFI3t13Qi/+TcZfdxRq9eYXJMk74
qxEEWyT/iPuNSoACHiPN3KO1eC53XadcfWC8xVSVJG6jwYfpQjUSMAEfEtRb4G6g7OxJKBevK3MQ
v4/EozH/4DA32ogmlrKOw4l5E4XvRi/aSMxUGFRSsI882VNvmdiVz/OiVR4um8qYdMnp6/ApH4Xv
dqSAHKUnDdwRbCupNxyzsEUL4GaD9bzjr9gFG13TfyozQ2k0Ticj/PNfNVTcKLaM5imfWgXIbvaU
8TGPtgF7Ouz1+Y75YGRdF8iPbBRMEUbqNgt+NMozXpYBWnEYX14RPAZmL6k75mryFzkgOXTgRYzm
J45h0EuV8FBk/vEo23ma5BkJ332PLVw4R47GMBLAuKx/oynJOH4Wc1aI5hZack2vGD74erER8EZu
xuwMcGElmeOtVKsV1YYOcM4TwLrXGBBQu8tJsjq3DwqAB564jm8eDbNCkNMCsjeOb+iJe4TPzLlb
WdVqKsYw6BZFCNAgfQQLa+SPAvbakBuLqt8RjsIKhEUC0piaX/zIex2+eac6QXc5/YTVRwRb723C
f4F7b/hxbNDVhSJ/sLTufw6QBAw3nPSAS2LJEa+rK4eJR1lABr5E+4NYRdzHb+1BJjCMsHUgfTM8
HkzoPpXXEQdGtL3XRsh7WHannK51tboKxP0SJqQQ+xzBPfwn2GyP5uIkGn+rz3kzzQleN2k3xIl5
wELa5p4zwZwWafVPTSxSMLfqPbVxb88StGN+dYErmvcCbuZfi/8F5LHczqdUtT4cEd9tz2BOCRMu
+RRAwFRdwL4mmyjScnUGwkZpICJL+sxbOsp5KtCArHL/WxeZVRA+thm3JAoTjHcEtZOWSk5N9q3p
piBrYXxgV8L+lRALPfWFaSVaHrpMxoIntu8dEEwDetQiRteq71lihrjYD8v3wAjFedJgwukUUF3y
n+3j+PaD+Bbslp2n3q8rmLbAO2jztrwdRLKPD+GuUJFn5AuCmv3MINZ0FxXets2OgebzQdqA4+BW
uY78mG6SfMwLxKjrD9B5MzoFvlwQrF3WzpKrhQD0gdNorJcUDBkPBbaQpC0cyW/79ptIMTP/HvzM
GMdbByU5UjRl0b16ajmB9UZet+7jTPx8itQibSr5JwQ0qaetXypKYRCWZPlUT4dcNzFFfvRO8E3p
4XMA8rEQP8WttP1GagSUFs9H4BUMo+S6Y6N2492zPRj/IPGKvsdQKvInj3t1eXAWu8gbgTsnqe/L
9fGFXzi0kfFH0WjZjrardDWEGxJNhvzaEV2k5GjCQTS2jqY7EpelK9q87/u6v0yDT1L38HsBqbQN
tmwtQFJLhJ3FadPQ8rF3Z1C7fQEgKgVTlvL8Nks4+bbKM6U/oqi1lG7lDrXSae8iAEzbq0fAFWqd
twFt6ptwFz+HU96YMcG5MxBmK2mf/XsrDKWl5cGyl0l5MpBwGvlbBMxH5jW25vqmwQimwe3dM/uj
U5XkL0HHIWojmMFtNHtin5pfNaTdCt4XyjRxWQ8TAGI1hgt4BFEN3Pa8XUl2SXJPdmZ//O4eXNtq
EBadoQPwag2Lsf0r9YOLmJj9WSwpkv1v/unf5rZx7cBcL8ZEFIqFqn2sjCX8NYYeP3ofhClYg1Bt
q3cV08l1HE31/R4xgnvHun9ySwtcwdLi5izZmwIfYJlczEHvkmjaEE9rbpiwKdsFNl3IDZLrLCHq
DeXsJJDcV564w4JTpr0l/fm7LyebpIsCSsAzni+ukUJYlAZBBrTL3tY16PRoLgQ46DgjXS8qjsid
1jOq+1kGmz0zEKJU6L0E2kGNUDjuRPnJ3BNLzVEr6Jbj6Ecw9eLy0I01mBOl3rlrM7Z7Q/5bFfdg
r8j+dDazITkfLR3TMNHP5jVu4oFrjYLi2IQl0ufBumIs2RBx1hPMALHjxyPDN9YhtxH8r8pwxP5y
A8IXui91UbwGy4qaud2nN0wHc4Az4omeIZopYpkuAq7ORHrhclmAu9ZiabySCM4+mHoh48Glufed
0AEp6SBYViMDiOM9JkRGKMzshpqjhVqgVHH1o0V7fNSwARLj+sPxHMMPvp+kXobbt3jXnTGPoPmx
G/opngPL/NgComoUF85i3W+TjLULLIszGYlbRCeMozfcNJTllGC1kG3TS5+et0hpCXwCKtocM0vO
C1XATEfavwckhthq6EJSVrAIynHTZHosU5whO9zJvQGAWlpDqDjErjsr2VjgdxWegyPB4DI9jYkP
LmQN3eH6YFJCcWzEqRXyKwGWhe78Jtrrr2G3h6yYR5hlwghRXNlaVYuPOcYpl1bkOIe46VAVwNTA
xSz/7eb1xK5eKd7xkHTYxrNigK/bqjb3+w1twcZag1uqXq3NJ2Wx4e+etqheyFS6D11TbIkYjSPY
tIyWXZCvulGzWZrAR7n9JTJlSZoyNWVFoEsUj6k1OU2KLVbO9GUw/+FucrqbEBXR+ew5988iPVmx
fyHy+p59LsM1dwvd5WfvhAwcQ+pVevsJwe69Fs/c8fBHTizqcI6I5hwzmqRQnUiRXwV8G35GGPn/
SEuiUW7X72yAZ+sUkUHUUOjfaOw3Xok33K6eccEtwsepy4BmqfiirbG8vMRN0oIfGXITvWhasOPJ
UWcL+UttfCAxHFouZnkaoyByjWDl+h8TKAfAi0pSRpkoTUl/JDyxRWaaPieSztFovEplsEzdphtY
VcJa0H1go2/KPbcUoSvRmajk5C+usQMxdaW5xe9DUwaNHrSJrSME+NH+1q6jrGKHARDZ/CiFjbN5
Vcg8p8idDtw8a5MPczws8YJT/pjXMpPiXma2saen8aOjK9JdCRHOG1jBMF1UTdxM/Ip5rbnO2nPM
NsfJ+0gsw+vXSOXAUTD9rM+vUlAA94BF6wk+5yaT2I7SLDnzylYP9F2ENSsDqFyCnCzbVuQX6i0q
44x9aCrsXaOoNWju8saWW4n6NGH0gevuSSNY1gPwetFRX2MLP3k3zx+JXQv5cv2qObTET8saxeSC
wweFnneIkNwVoG7ajpsqr6Xeok2wHxzabMTkYdbeDx6GBmDNvnL3qasCRiEXYA64H+ILIt7Jun4L
wM0x4gRFT+qFxtxydB2rA8p2M2RLY7lx0ZFUaCWGg0SHfewkmysvsNEFiL3Z8X1HkE4kM608z8Nw
ZcfL8wg/qU/A02cTnjPwyW4ZDWgWPd7D7Qi/B/aXdfzL0U37Beq90RtyTbPJpqR8PHoWd12FzOR+
HZ+e117rp/aRsLEkKbiBjwCEvSomhHnGDKoGvas9AaDFPEHHTmb/fipXUj5LUaQgAkNCbs0r9RTE
qP/FKhFmVD7zhojTz5GmpM4IQI/rZY1KDM9Qx4maAYUutsQoMDEjKGBWHt0YV5kWZpWzBw4jaenh
mbsTs9/X7pNXxUrKvaSir4kgKUmdYzYvAb9J4JISRNSnIc143Ct2aWVYd8QiZnUO2eJy1VLdZNiG
6k/RAqTAqE16Q8nvwLOGkTN3QbdHCE0mKboIwgzz5MNwaULG8NdX6ZmI1sEDbP824qFPRLD6DOxj
w+OZKiX43AbLHReXv9G8zw+cp6MTycy+CNQ5Y/IewQdxuRHPOMzFjFA4z2Dkh0N8+eMaX+p8u7vg
ntvVac7h3DJgsz8mDgZk9FmUXf9l+Q/7XzbsWaFixU8XKezEpPsRkHov9hJzGH0qtoi8PNG+SmcX
tWXp5tndQ543VFE8ga71xyz/8e5wvQzdgYOURnQph+XmhsJrGJn+d7UyNHE4IwR6VwSFSErgr7qz
y6pqnxoEtIaYqQ9AmPTMgWnPnDOuAgK+dFD/Ve/h9a+bAatkUWd/jchuNUqmnEvi06+uVfUDQtIG
DbvXyJFKIYdLTxfu50MATh7DgioQXJYZL5sGd+yZ8/2JwFtA9QAKgVuStbx+U89uRLne0103nm/L
zGAmzarKxeW76YWlB/WYO9OvlEmcfLqsx2dkhGkgP0l55pTwg0zt/vzZwOye/Xbd+01P+w0pwsZD
SdcUkGYInFEvrwxK6r+PHUusKU1GNLCaLPs5aTb0WyI3w6stsOf3/0WxmKF0YSbmXL3JQscp9zXv
S/wbYaQD1AreEMQPWRnuLRyZo8voE5m99E/YkEei3s2Hrd6oL+GFFECSwsPaN6tUW1WeIZhhu4NT
MBF1xFqd/3milXT2mQMTsR7m6KqJW8stlvtJHHZ12lzPgy0ZvO0YDx/q0Zj51icR8fleNLVh4FBW
EeHjOKmaAy1cFMB04YYMEKbzCFkEHum7PiHYomx1IzzJTYwHqHE2eBFRi+qWXHoI5cQoZkqoUMiP
5JoOBnpt2ngQumJ15uv+KdtJ3+LwtR7xDk8HG2GwWSUJbteKLIm8HouzHl/jAfBN/fFSW6yXqvuV
lepRL3zl66ciwIt6Q6zz8tqzZfbalx6erydtOzNz29SwQO+UzMhT0hS8I+okeWelBpTmajKu+jNh
QRD6mcfR3q5UDCzZ/3KSK2/cfkw5KuxWYpU61RQo7WSs+RS11wkkJGJy4Qf+mF7zE9XxnrpuO2pv
7rqpgRBDhFnNybawJhLL9sExo2gJKkAU0l+pXcgFKguO0XKwbatveEsItAhCARg6X+9VhwEnimF1
4nt+OE1HSafMrqqV7bJrxbTWY2dBMYDOoaQdImImo5zg4+hZZh8nhB4+38KsOmY3leF9MkQiqNyY
WpvivV9m6uVuCuBAvo0NEyFcV+IqBR5gRFR/wFChOjqkE7G7L1W0mjh/ud+vDiMuKauL5HyiFWOn
YxBT4XPxDYNmvd3XIL6U2QzhQSLo+3AZYzS+/OJk5dHJE8SeiJOP9iVTmHn3bEcdJ07oZi77Pv/g
it1fnHvnxpCFAyXTYFMyZf6pnqFhOSQv+X2VDE1p7fY/7448u25OiT6++a5Pm/w0RQzScSb66iwZ
B7ZwYLF6ZYugtd6rLBBUGz2Kqq2IXkPVRRtFElCPRDomuClumaSiAB8eonkOcSZmOIk4aSybVo7V
jxls0zLPDr9hZqLNm2wZS1qrEevnKrWzlnj1nrWv4Xve2ELzF/6xsocbfi2F7pvhVHNhmpYzuW3a
4z5RwUo3sUJ4W/TLy7vIcaJaoEO87iW8p2XguwEYHaRlF3cdsxWPZmh9/uyhhg5I4ouShb3K910y
iByxVjjBOAVCEYPTgV4ic9LDf3DcbmfFqpksXxlEPOEo4LQ6UEjdFf3cgtX89ijABp3MBSBJnJmS
ZlDwSDPOpTqFDceh+gxGxmm2/ga7fnFH6nbSCTgq/bsIqg/2oA8XqsBXnd3kIQRG3g/owGK47aWi
04ujTlRDnhIEU9efa2iSryUXoMUBOBIlOmq6KFVjvU+ozG7dbcH6EOhnQSZKnl18BU0oiUKCZ2Up
fHB4ko/TyfGPi9xAkRDSScbQpmW+h5/C2Ml/kZdPG8T+ERFnCkSPlfcMjh6RX5MddCdtdF1S7tnp
ykLXTAopSi8Ldzx6NpCovCS0xA3jK7ddK3Ols0hgAyLAxlR0cwsy+/DHZrTavMnuWdkPoDtdh2uk
brHrwJ7dUoqd5zQVOtjgn4gsTT4sg8mvBz/KBGZ3LOARt41s86gXKMfphlpov5/HTvW8K3SEFU9E
O/y5oy1hjLvmis+VAXW9GQgoZRCPn0cbZGMzeCo6UERke4AnxCrRHWtP/LFt6aTq4nRIoOApxN/6
LRu5/FGjTxuRAc+HrWn1cpBLf5YvmyCfOX59D24TO8Vu+rrMMO61rsbZgV1m2XxMkUK4GYb4KCH/
3dhdG4AGFysnxDCJjsREhBDVvMH+D34AVcLxcgldGqEhIzMxA1jMqs/zcXNY+6mkXxkBzUBakSYg
AOIkrsZxpfUUF8scOGjcNc4HUTKN4zxOs5bN9oePZqE2dqcm3GPT7aecaOGfcrBsOJKn1TEtik7S
9BnVlBAW028oRmtpOqggzsVsB2my5Tl6bo6O5Y7RfdbmuloQb5q95CeM71i92rTgOAMv7BVDHmef
1XaHlZMRQD4NpJRfDCuiKa4oU0Buigl5d4bjZOQ8IHp+zbtDbSGBHO61ewwwf2fZbiAVSwG1NSgW
FCn7IpoDOfA6g17/pZnAr9R9PsU8kWvyR4PSyq+Y6GyQatJ4GJeChxn4DnEWMHITiZvF4wKvryNX
yxFXaBp+DsMqwRsAlvlXs5Uqx0afCJvZBbT0b7mD5hdWvKZuNoHK/ammlhW/YOhV6vnZQaFX+8jO
eX32Bpa1gkG6Atu7VgBI6ug+nW40ZZIDzUTXTGwB5tZDVV78TZvbXtskMINMRALnqDtr63Oniiyf
fbI/+6fAjo3OImCRb9LPbwbQMxujBWeYcPi/hfVZF6kFWWLdkkK33q1h4w294kap6nodwpSz9SEM
CqCuanRel+PER4IvDQH/UIgJkibKT6fZot0TJGbv9RX9pgrUcw6sab6B8VYM1+blsxPq2tRsOl5r
UaWQ0zkj8xID0jtoApEZHOmJD3vqIQB3jJGJ0OzkqQFfvEbWqjGTfiXIP5GbFTS+9YgMPMopK7Jq
S0Lh/BRyCaOEJtCTnouujcu97GqCSlpC3etJKgINGhQyR51EjGGRKmc+3MPaih+6sXjpYGdyn8Bw
a5qG9Smh+ZGdhy4qbcPGwGFa8k3hQ+N2Qfb/C0NXifQtkRwXZu7sQcNIqH7GWYzl+AkJI2B/VDEG
udCbYhyPQNbDKwcb48h+O4OHSBC/GhHoj6+/n+tecA3LKDhDK79o/BXkDftk/AoJLniB2zHYzNsQ
mdNZKICB63UWBkO+98ny8onUkDz8LPGbUBxWAK/fa39ThOIYbP2nFub29VU7wtQD8az/4Cb9pser
LTlHamUsRZdmwxVoP6K7641P30wr3IVtKq4pBRcg933blyS7eD1HhUSyQOJZfkMIAoIYWfczz9gv
cWi9pdL9G0qF2d9HeZ/Xh+L7a1Ui5SWDRErXPzYyTGbvyrkZ35xYbhbFxqd7jcMi3URHBUlqDIAI
VGZGnssQmHqC531GVxafE3iw0j+4XatOz7WY/XIwx3LkhMfav8QmXWmN4Pf8gOyFZqw1eJnJXV/n
2/WmbljiYJpI4NhS6vQp1d8yNsvo7L990Ze5fMkKZfqaDSB8GP0tKHuLm16f420sPHL4XqoHganW
mpC3C/j7+FB0fVHgNk2yu3rH6XpdGzpPuyd4Ste1uURaljDRktyzExdnCsyb5nb9/B+tcX7gKBDh
dGczZ3xdUzkSN9crjhN+E+LqP2ksGwQX18LLjPI9qjmsU7Go5/ti5SgrAucFrcoZgu8Jy+SZV0Eu
uQ92vqEQ+mrWqZv6c179eVuYa+NVSjqwrwcwKf7thM0QRhy1lJpG1myjyxsQIFVIt84PmReV3LV7
pttvO/e4BpG58HW1k4vBduv+4Snh2wxbcpHymydeZZaO+UXjHxm5IrYYDjotq+31t1xM91p6JAjl
oLHmoDnEcXnvwaYc/Rv/VLmpXztDYSHZ3Yyy2y5Z6Nev9NbveNwfAEouIyxoiHCSSCfbSDcxHi4Q
Ejibu9yBahNaRKtg4PknH6m7KxU+psU+8+A1p6CFSgzRMksopaAAw6M8evBzQnAHFdebR0v03Ht0
Uo2f9QeWC3sou0Sk+94aHcPzcXHLxw1KKrziTPLfICQd+o8YVfqjEvB3OHFlRT4KoSiN0P/ZLESv
B9uHtIDzT5FnX+8Bi5qagLLbXZY3Tb3ETWugmR2rjRADsDRz8h3l18apO+uG1y+BdYsoQT8jhv7i
P7yrRuGMKJCGXDjOhBbS5VQFeK2Ftwc/L8+YzPgTq5DczFgW7SePcGY0u6TW5j5SuaEIDFFAHsVN
4lhnZONXV45+Hcb8KarPDmCdgfDrbFcQaORgdKEtXYJsXwit3BdaSXzXxUKCCrs+SkgXNAH9pO5W
lxXm+/NU2NBnUZKoMw6SFB1EfHGhNcnSwH/LrNQrqy0IU0FPCaCsB8hu43t2ayDi8/we5KDBRMpd
/OTLcE3MncYGCS7lyQXltz94n4y6xMkPnhTrZlZ3ncmw6IQGVjRJkKrZxlfD/k/umflzVplXaRvT
n+JzrwQ/RLnvR4f7pkD259KARFo6l40gQQ8sCqRuYmDBKh/BEQIRgBsxXPLkRSGH3rpLjAqFcGGH
OU8orv8C29cvL/5vLAtaMiIwXHBBCUY1VQXAXSfisY1YB6lAFgSAdNhu9OSYvYzgJmjnGuCXPsWu
1TctN19j19YLPT+UflVvN3QjNzMZAV5iH9bDYh9+n4Mazt7yTTKj2g8gG/tyHVpZKlp5vaeK6HHd
rGBX9k8ysSP6Un0ppG+sRe+zAKrIRzTmqyHxFvL238I7X9Ou/sCzh93tlbe5C/CQ5+xXFez8EA+Q
p7xDXLVtqG2kLtlivTNYRqLyjK7YU+X3UL1PeRGDPH0FhZbG4smxkrQWcUgmyA0osd8Xf3fsr121
s6+gw3aXipxxWSjYnvKgXcato28yoaZ7zbI+5zLP0YJSWDXo3lo3vsa4fAiK+7nx0Ig0Ez0/hx1H
lUGvF1OSKzD9ye71hNYMoUrJXqGCfcX3xf082HXrEkht4riab82yM5HEtLXH+IO3HzWcIWYiYqqb
XlF52/sc02dZHcl7DkHpKRN9SzekqQDUpVYgFSOPswWK7C4/qPRO9QrbplYU01JaJbn31DQPKDk5
FTnytON8riP7A/dz0AGTjPbVbix+KdCb2OTh15hGu9XiiWIkGvfU1hnP9q7pw2cCJXW4baqn4F/f
4sbvFBH7RfyRXclO76+tKTu/GJNDU88MSRIbnANgnU98Y67q52tzjvgsv0u+75UtvgP0zTltMKxb
Gwl1XvrVY7DItBFgIHfqfReGPINgPJXbQdu0k5pFrKdKs94zpwk/UDjIqeLNpVhiwSiqa7NH73bK
FubBnNsiqOjyDGffFskp1Z6Ror5KSbzfrqyXoyPaCG4uw4wKbXDw7kZfPCwpd+IoETun0HQI/xX9
xKQ3kDFfkcSg273mYfyWdfZE7H4OHGMQ2+HZ8bVSydfpylQD+8TYixkRqfq9X1n1evz3uHi2AUIV
eALNcKkQdtPlekhv36mP8tjmU1yLpwXYxGxrYvQqiGKqc2h8iUg7+pL2zb1ewJ9Qs0P8X2MiVUHd
2Y3fqL4DwQudNgRDK72frhVFlK3VWkTTp2mzJbTUnUAjZEuzoOZJ6J6/jKj78FyQfSu4nui0Bbt2
/Bd/Ga1Z1RZxDx4iM9mbOVez5dkjhjaImZK6fOlEuST2K8LlNfZ1T/2rpqchDfey+r2VkqMyQb7E
aSOy/HKwfbQDfq2EOrid+bnD8mHmv30f38Wpw/fa+wS0rO9J4ojSv1KEaabO0Uur1CIpkVkSZBB0
y5vmosxIR4RNivVGmAPfdSgBISa52agdtw0F0jNq6sLpUwFELsrS6pa7kTf9CoqbuUfrlj8+Fe6e
TBxl0TxhhwlPy1EkHjo0ejK3RG58kLbzQyB5ryxGzkzC9xHISp4F9WhIz+vikYFddAlFKBPYs3vT
+3mIYGahlRa8KqoEDbYRLdcED35WpRj5X9/RJxVlIWPSiGeCTWfndHDS8VNM5oDL3zRPLlIcIlXJ
TdxSGHOCQwkozLJkUdjB5K+WOkvzqbMPKIqwW/YMEbDlWbsIsq8OuzhJAH6xHjddfTx02EH5i73K
KnGAaOEIAXmuKuTYBiq3LDgVMFjigmxKKPpXYlRHjBketP/PSxtTaqFoFJpVUko5eM4JBar7nvOg
DHQJWM1go2ObN2XWgXbILSxmVJdSb0CSju0IZHb+VtqG9ePuhaNcemccWgMgwC3aFNqCRkdz3KVI
80cLeCwaGI8sIq7tewY4ICEVhl65oa3LdCAfUvMr38/88XJ1WFVFkdGjtpNmk8C4dv7+TW4qiBcQ
nPHInb7MB1bp51pvBkGFlBYRIboD79fU7N7lshjo5lsV+ply2ori4dlKcUNvMsovBcDuPPT16D7+
9TPwdf90/xCl0yvqATXCgtspNWbVLVJlKAKLJ/in9wFmwBNgr9Yys8kGCBU4C/PRbnW+B5mSvDOK
qleXbu126uZbupRCHOdt3r7WYDmQrl7NqmVzs6b7MYAEZtXH5NGUExYBK3SLS3acQZ2Vde7T97QK
/g+ib2XMUcFwRVRWgV+AQLY+J6JUQMXvphg+tiAvNNgaF7CtXmblqOvTAt+/4yL6iwkoFlbdqVeq
ge7sG0duY0pY0OaknvddL717dbF28PlhPBVQtawLoMDjyzp0Cka7t5c6m+X/WFjtdihuleEnglom
ODuQHyhww6tWiNkHezb57/NpiUyZprDcpM4Hc6QcE+nSmFFGuuKNgKUNdBjKuFb4DqAyIf+G26DJ
t553kMXoDhxi4IPbx4EIRjEdpN3WQaZjvqAZkzuYiNaIKBN6uYU4k2YPdGI/l2kPMXEfOHbk2dpG
1vtdjPsuet7IZdbi55JAedP/LQaPtzXrnzD0D3Uq73z9s5dBz1BGSKzEyoDaasYMQH7AzDykoQc/
COwCo3u6ENVv26cQtwGyv1S4QLa3t/CEQH8EYRe9Z9Uam8KFK6qfRZv+7Qxu/dHDTMKTU3QrkDyn
hW6Us2ZnwbyucJbrim9BJVnZzzmpJelJilUbyS0K+E1MCE7HmtCHawN17LAIz4Ds0+oAwscLKAXh
tqzrg7SBQeD6/bY6uh3om0aLVNOajrhRjZcZHxdvfCRv2nMHLIhSJF2S22BkFGWeyB7L3gk6xf7I
Eg6j6VBXQNXKsZljDC5Shje0t5ZUTctAuWNNSS1s29CtAfWD3en8mMxf7G8xHCdMEMQWe6trbJPn
03EiCUosPnSKlZ+NRJ8MPmr3n8LF6KOP8xzy1ceQ7OLj3n0K8xd9T0/38F1I5L501tGvOFRGLC1W
c66g8U1hxgqh5utIhN7neSTGEMqfk7ISxL6SbmppKwLDVsLDDBF0Sk94rnOO2OhfqKA40I9Kee2i
LjAYkr4s10/xl7XVbtULncxWdQg3UOJsXVkQHrjIGKsqRpmW9gKkOCeRRzZ3xKqIfL4pTU9oLtoE
4aCcLyqED+8UuvIy+2/PcDG+IHs5+oL4RhZeL7PmCSilYDkmuQew6h1yfGNVcbPk37EuKTELDBoL
Xv/D9ph6vipZfFMpnY9r0HXPHkjEssRFFdwmPCkX379P/HYeC1FnpO64JCYdjhHMIrSvlLNnwSmz
+MrvKJAX4uM8iSbQKjMxK7PamXpO4pU31mkkWq0ue4DR3qiYOKIFemF8vCyTle1BDKHhm0kqD6g/
TJvMyvnuI3j3OyUv6LOeTEssuXAe3jtcCN43z8V+0OjL5O2RUjdXJhb4uH09LR1F/HjXSQrYvCVX
v0Ok/hfGcsKpBvyPTHGolnGpJ6Z3yFHcUiXTT+DwjXM8+CkctoRh9EJ3u5J8DYsomgmkTXlqEeeP
7xRKiSyflrl33QWUah4co91A50f2a+sSnbKn0aWEbDLz6JlGQzzwsBSxF1QExx3f5KYrgETr7PRC
zpWkKIwIi99KbjzdVgsEer6oHbbave2yhr65YaXcwQ2BYToKb9Obv5KSWhgupvrFc90THu3Hzn3X
DPGTZiSYgNxAklplnnWv7oqNj1wvvDJyCqCp32o2kFAYyxnX+l97PZ01+Rg+r6OY3J/MMGwX9Pe4
zt+OvEYyl0MCmRtNuxCdQy4Oz2liYWbvOHbleIA/q9tQizcHToNP2TXwWLPUk0KltsiCG6vuF79y
VzpNKqEO0fWTp5qiEYlNcQbCB2U25RHuexB7EKTjVqvGCnRWe4uzYS7wAHMvNz6eCpjmRwveGIqt
RtE2qT9sSIsYjH2W3jwVLD6pibbztvDsRRN3Y0Iw44MnLXEk/NZ0kZaD339PdhWFXw11grziIUZk
+f2OrylarnBFq4Yl0JYjO5WF89fey9RLXcLpjpt1e1EFm3iHFDHDEUM//ltBtG7UIl4UmYpy+hVY
FkWHNg9tCll6fUxw/J8iklkh66rMipzXUkL0BBzr67Ap9ZEym6qmlf30COM4QG+xET8ntqkf2etT
/+CTqM6WodNxFCBcNFKCB7FA9JHOOh/m8Ys9EMXAe6F1Ky89LlJicufCCeyBfUZIl/sHQrRylOtU
ZwwZR9xOp/Xe2m/uzCNy/GsnI7XEx7ufuaiKvc9+UgUPN7vgQhPUSvJ0eYLRX1RPfqOtmLKmAv55
u8x7I4SuUUiIhcPFRZa2KCk7kYAB3twIA2qcikfRpfFCtdhatmD2RIsypp2Uz/J8IJliV12R0A/y
mCCOExINpwj6a1VHnvxLkIJgHqbBi8EEUgjZZPR1vIHhao6aHU7g+IyVFCAZEnwKB2uLIb+R0HRl
82qAUhdmvOcJ/iFyi0dH95gMYmwa2GQxMjiJFqKKc3jmaodZKQyK7Tv+cnhushFAzOOPAIFAzccs
4Fc4NfAuhJgJfD5htn8+LrqvwpoKdOXCUtzns4Y3NKpFDIQHBGzMd/uLaiYomUex1KGvkH7KX7W3
pB/55M2W+1rOv2UysDkN72PK/bi9AP9YT2WagxAYktMjH7mZIbkDmfr/BZ2CpXHm246q/S5DXY8j
qHhWjL8velWRb+plxT6+q3N5NuHF7zB0shVtW1q1tkItpRw8+MpYyXOxwA1bPr/9ve56J6+KNDNi
xl89aabiAEkv3Nbn+Xa02Mw61WlNOEa+s+wmjahPR9HhHN8x3yGSS1VhO9Dkz3vzg1uVaZOIDLUV
LwgYMm2OPs66kGM2/09ZNOAQH9dFWr6KuazuUi3RTS+MA9M/OZaDi7h7ZBgH3/roR0imTnQChID4
v/nxpwDqKB2wUl9mUU8FqfMP7PaPdnrqRIVMObkXuHTdZsvVCjP2TzVxvy5xclnqimY1Ajuu8Lhg
nlRszLVfPFUnZ5EuEL6qjSYG+1x5gv0/8+jidnkAevhVVCaIg5/9l3OEbZxuTHEhbRk0FXwyPSDt
CE3x4zhfMPY5hKhlY8vPUidd/g7cE0nEKy+CqFZgXmjB1iDrl+Z8tduj707y1ExBTsm3pQcjJzKf
pTR3LQV5TJLpxSK5TVTi/K+CnxT482z52tdMpcOwDLqRkxQgHpD9bL/QzXdybfaPNEyKOv1ES4gD
iotpfjE14QBiHGogXlYgaIoxvW4hodfKeCeo67BrZtPb5JBN8sWylswwV0PsOW5PlaHiEpcDUlkt
Ky89t0J+NEqnJbEDXvJN28bOwh/Q7SyPKWNYJQ7O8vAtW1HKECQTJtH3pN1YW2bSCmz/jJ7cNXGv
kVaOhF9ud/MmeUyVx0P95dfH+gCxzBusA9ntN/mVwbI5OcPaWIAFDbKERba2TxcLZW2xKJvpFmYm
VUPFNrI0LEouwFbnxzmTdBHZDXxnIw3UuMNPbrdJPaoQSoFFZByf9eETMs3LGtMeSRZVB/LRnWwK
3nHPRtekr0XxDHGgRj8VqWT4sAgUhWZlhtzH+h7xqJ7LIAaKVdezBXlxV0VvnMbWY7dM8UlmyVvC
wBnc0tt7atpDkwgZZLQiZrDRKk9Ouoa546Ur5QXXbCM929CtIw8Z1YckXeDg05PmgiiyWPxJiLg7
bjHdlzuXRLZmbVFPfX++/hsLxiHmYGLIndX9OKKzPysm9gpag9xiq+jTgfnCgLecibnK0qIYvnmt
JcgQH/xavIjmojfdl55ITwlPQHmMhPIu/34O1i6ps9GsdkeN8zZniC6mL43Gq3Xsp3nZGrb4WMVS
NOMzx7qV9dTBcFZKkDMYppa4kGTWvQ+S008H+nYUI1l0Qr5gITcu0ZqgFEzAah9O6BPR7UAva/f7
B4WXlXUiROGhuQzqEcD5Skn9fwqK8dBwMxx8xpvm1thqIReOPoLO+tgsuAr40jtxfejXeuPXbIFc
njagFLEPhDYtbMecH0yscdLUEAV4gE69s9eSAlTuZOsSowg/ko0y9fcJcmHt2rqpPBaX6hJ7hFk5
Kw2aQeH7vJHF6rGV/UWJ0Bk02rTWHvDK+ug/ByE10F4av020N9LkWmcjbCQXroVgPpolrcIUbgBq
PD+GJvFyocvN0oxxfqs4zJtpqOy7dQP6foodumdJrTRCQxwuqFPEEMCDhK5up7Y/qfr9uK+n6Z/x
E4EN7nvE2F5EjCtzF6QsZNhfszrnYORXIbRiyhCIdZtk0Qju7f8pSR4tmuTHYQvEtrKqf2Ms5nks
2mW972qYn5t5/4Qomg54Jv/VLrip+xkC99QuJ1zo65LHrX6dpqq+75Q2cvZ6XQ8v5FePq0lF9dsG
BudzUFJoilwPNQHCGOL4jZagMUmR74cd1E0JYQHUAjP8YYlBVkrMJURUR+luIdFnoUD0HFIMZwEw
PG1ENdOjZa0xfRspptff7QyXM9j34HprQBti81m22l0PQk4k1jRdbWErPKv6PS9k37c2aDME/pL3
M+P/jy5ng8aTQyFo12DiVP76G+CitUaokwB9Swn39f2G4At3hq4vYvbeVCIKh+VQwaQ9WJr4SEy9
SDrv8/WScsU+hoW0OcS8+niX9ZcCVEFYrVpSavr6/66QEeLWY3UwUBOg6XEUNYgniabtiCoeF5IU
+mB62vhEuvW/0odl5aMjp0NZe4bsOqg8h9q/OF4hix0Usy3JJGeGstX9yJ8yWdG5UyG4csEwo1Eb
KW9Tu/tsXu7+vqDfvW2enZonh/+gN5vefRpVcJHXJo7Vf4qJbQQwKIpI2ZuSn3pfKlCmuJESkF3j
/FxOi1Amyl0afiIokLdtGEeRiQyR86cfEq1iFRgLah8lgTS5CLUQraLpn5796pB3/okrUl7hAorq
uo7eyPQp9S9CxB9h1o3Acfkt8HC9DZBHsvYJkR9VnYkGjAdtKymiPMGC1+/jn/SK67ffYcGbxjzy
xHwxIJTZNTyX2YZWHUQ2/ARjVpxUY3i0ywzQN+QzWVIsMpdje2+EM+b9IVhxxNzxfGWj6yPfrvET
2DewlfF3rQyYZn1epaaRGDbF36HNkWugMV83RaDrC1uVpJF0pOfHfIDsaiih3/9YbUPoFhs2o84p
PSkbjwZ1Riwp2/3dslIUda/2Nl/8RAELNtFDQ5z55l5CaiwS3j+OJ0KrPjml12EBA87kdw/tBUGS
AhZKF/TzGA3xn99HIjstr3klLPvCq34IIYBwUowPgpuqJc8vxyq4t0p6TaltkVe5INEYkYBy3bRZ
9xzinVi6I04XDt8nOrTvdwkGEBe2U7wuvpFJufsbWZEDyOe8tjgrojeLnQqFPFtpu2uWYrxDLnwZ
d3GR13Ci1a6pEnda2rOMWb2Yh1eho+Ee1DpMQiI70biJeuLvs0u15RgsdmtNoVfyNJJqWncUzZYt
hyl+XZe7cSJQieyT1rn9jI2Ix2DJuFHLFgaJUbbIY0Xm4pG4JHYSi07sFXTFnCPYWOcDm7kqA+jD
vRTd+cYUsRE8E9gOgI1mbWoOD4p1Wq5vyx1mVZNTTiI5lzemqgc/T7ypS4fK8zl5DW+Qu0MCCAgj
6Q/5OPVGR6vY/m6CjS+2yB2IBH6pumnKA8OD58R9MWNMzy93A6pDZmAMo6xNAVuqDz3XKx6c7rZD
Ey4XIpfHY7BQ82j79bORT3Sx6c32dM6RWdCR0Xw7yL26pnmlGn8c2R9f4727zdbAAZdyQg0JNVDY
nmrAn1MJyz/ftd+5dDDxPHAasShOThzWTpQh7BZR7GWkJsYPJ3AUbmJ4RG1JKxVbwPx7BRHUqwKj
TDcLILLpbtGMXtFT87Nt4GyskB7FwfYGcM9R89uqs+xSLel7mGyFWG6KQ4D//0PEVN8TuziUkwA3
o38dzSf3FEv6p+uMQcMqQcKbi45ooze82LKYzom6n2Nn2VLNGk8wVOeOzOj92JuUdaGpqVxlMgBr
MyxRxHBkLLMJzSvj17UQbGarNUovbmxdSNkrelX+D+UmONvGhsJger/F90guakrI11mzRCvDMGXB
jZDmjcAnb8AKjL5uJGjkRJ8JxQdSlSUBz4qy6I5R0EsYok6huvjVpGPjmlB62vI+FPnF8oD/wVZO
zBO1NFRRm5fhMegleLdU/ZGFialwRGRB7MAgBielMWs0U5vPEOJwAW75sXNTpbg+I/iaG1/sTHZC
7VVT5JAP3B+qbEw//tEQ4lbG5TeveOs+EOU1twHV6UR1xMd/qzrQfKjVCg1oo1SzmcRs7TlazyJW
24lFsLYE01LKU/rM9FawEn6T63lkIxk3GdwchbvesjLCwzj8GzWGAjBU5m782gyjJw9g2xLnWid0
hHEaT9YXS9Gyc7XuPr/2gU5hPVSGJLFtPtLDaAWPdr+5nUdrJTcsIyxSo2ckWmV8KcNOLgpObv61
i11NJx/RGBj1/3txdj0q6mHR6A6UinFCak5/awa9vY4GlGDHZnJAxeWbPOMRsr4PGlE0A15TnZed
b4fvNpZsnNbhvf5JLeQ+37/9N/ULn/ie0UAiP8p2zOq9oCe3hwG9B3nOD9pn2eCRW37HO9dokcqh
SF+sStS0mtYAZbB+jBKiiE/hdBO6RnoVKb4ZMFxdU3aHD8HnVz84LBAB1rAMwX8+YFSltzUzn7es
nJeUZ7e3Cx9N+GRXPb5yjQaYje38rTxQnr/KiNBEZ63ieCfsq07voMgypW1gs7e0Q4IIkXLHviEv
iD+Qc4+2lg0O9tX4DRU1932p20XfjgLsFv0sNc1Pxh0Rsk7YOJvY3baqBIv5He+WMSAsdbgDTciV
BXxa4/pqLpK9h/EqwdAkw8XegvMs1OlCCP3c44Ga5Fu34BtLxAsuWZ/wQIWKuVbzrzkMwA/mnYLE
ZTYvpgfL0JWS5lgkAgCBGdZticJv0Rq6lA7qSMcQjG5K5a2UR8qvsQvzcrpq+YZHvaY8Ygict//X
APTWBbcM8Gj141TeSGMpFkv/tMVWxazTgI64vc2Mg4yJ4Lyo0ZLmU+/KeadqbomYc9juy6DPR3SJ
l6B50/fVakyL0Bhfpkd8bGSTB3Rfl7JGkQfgtMyTKt7ac0Kuwks7R3BK43yeUvJz9FHUcR0Eo7IO
N/19OhO2e8GD/G1yLoTS4QDuymmvJLwUpXsBj5vTQ+HytTxD6nl5zqpM/EP1kBWyYos58aB/OCEp
xpEZT4+kgcaYOJXH6AbBnt65+ZOcmU5o5EActAzjhiU0fZ9Xk7kL6aOdwMzfmCx0f0S1AGoeXAa6
6h/RxlugGymDiZ7aZynMMNo5VaoriEvfC9YjMxd6O2POG6Yw6MTSJuSUy4AMe+sr1oyup9FAn/k6
xvtMZKgfOCCDotiOYYixlOF6+u0xb0WIJdEjPr1VuA40+8CfktVouK4wJwY4QfZE4fbJqi0T7y0v
qOe2D0AztWkJqR8nB/Dggq8WzeHY1a7wo/cwQnTuPZuOQBT/FQrGtt/djbwKx25ABKBQ9HnCxVCJ
bUrcNHfXYNQVIioWE2YcijNWK5iMbOwsIUVX0hZDXPPNFrMJvq6yMkzCyQFx5lt7iLFVXjGjSuv9
m1wGgaY/KslRlLYo57PUBFF3Nrf1mTniXoXJ1gKYArmSZF6RbJniTuJ8S3dxBvKN1xbjvI+CVM0C
V8z/PIyRI+qQj/byLy0p4KiD5I8GAb4pL06+y8a8m2XpcltjDyb/LWiR1XWJtzVit2kEj9+3xxBM
5cRn5bmiRKSfjFWn/mB8zZCFgJPUFJhgVrHlNXMe2ES1kU0p+5yZpKCqhuPg6a1N7ewGmJC6zjRw
AUPmMHTk14Nbb+p0Yq1eXRzvkwli20EFtyynQiQ27QB355Zm23klp4W6DNLggxqho0lW+/6Bu80/
5yy/heD3ICvKlrKuGDF3QtfBrAH9BMn5Ban9/xiEZ3zzQqUr0Y49VBgTezFcKGh3vRgnAZdT869m
90roeU36wZJc+z3thCrTHoKdxFL+L2h8kvNyhSwhxhooenup3AA+gvh9KKp9WExVewORiQFRopTn
vt9xLsriqndaJ2bfM6Fnv3onYfBUQbvtthaLEQDmg09rxVV9hcm3Gfccuth6Inxvreyle5DBtokz
hrJY3ROHlTccjNU6+61hLouCewD/HfAJf63TyjF7pk12Jnw1E0Vkq05NrJNX2YHvC5gVfPJuVTct
vHSmP6MBXfZQ+F8tohnlZ5JN98CH0LvoF1NE5lW6v8TB0aCEEahFpVFaOIwqUwvVUvcp3BRUw/wn
L4z0kQKJSf+stc8r6TT3BNw0b7KBX5MqeRyoUrD+3+oQFTjzMkqdL8wqzyvDlt4aJgSfC9+KKeST
YjT4bsdbjZ8j6kcm4E9Ldoh4MgSkyIcMdklLoCMmcDeDHtP027C6pNsW4nGPrs9tj62EcQ/VQGXX
3Mgbw7OEWfifBi2/EaHCKKPqcBSZB2q3XfAdK4cK9ZxkzUSq9LTbDJ84SFotpdKY/3VPe/+HihyB
eaf38E/hER5pJb6WFgdRtDcuplmpXm1C7kT8hlGjhszIlsTqud7a7Mp1+U4xuxizEwnq5kviG8dW
zOuyW5H2+8qC/vKdeWSlEi0O9FIvsA89uYGbXGO9ydpr2FI448AtgAlbXJvfdfGOMWK7LDHEFRLX
WuifiNzbOl7fx3RmhtoM5OgYpTURHIWU1hcDUaU2lNkHdr9j3gOzVBpBt0S4gy+BR6QHG0fEUPR4
yh4p1JQqGHZg94+UkNamsRUmyDVTQmji31aNOxFq8al5H4lKJbArp3LkuPpjTUmi5OmY3fk7ywYA
KqAAdeineZ7AM8+4TOfAjLb1BC1LPg/ppseyuMRBLfWLEUHBSnLVtgKQtbb1SjUsGiBe4kF3PBvy
er9WVlZFHaML6040GJM2VMuhDjMnSAm78h5l/6JZYp2u7ZOSoRf0li7R30tG+2MBKmIXo0h8hpWW
RLkG9gGHoZLJWPCHCPpaYUquo+DMqjJBHwemX6pdkyDURU1DolZCkj+34ziCnr7eFezBoZ44bSnA
nkns351PwAKsKSV5zqWiUBOjYWHZtVlBlSzlIja0LD880wgFV+zQw9MGmQ4nw1luWvYUQJGubTRa
a37juH9i0WNyP+33Ujzj8wXGHEgb3XADJpCQVUUi5E/fi8/mozxWYQwltQ9BGXFxJGycrz3StecV
Ayd9feu2VOhWfRyHuZw3tnO9fdgIvXF3jYLUJ9P3212wzQ4o2bpKN0icqp/70s8NZ87i4QAtOYY1
HelIG8LY7+OV6s9iO2pjUwkH8OcXRFydqpbjc24Dr/3byxymUZzzeMCMIfF0GbEz6SmyLNM9r/Ip
xvuimjbi0tNfOczBzsi4NZQk/TlulSAbMLNaaoQzszcQP6QbiKMy+Z7zTVDImfE2E0lGFoce3/Wz
i//1Uvz40iLOvXXMibpy2lAqIRA0tX2HCu4WQRQnCHW4rVFGgRB5ZcFqmAiLOJhsvApo+0DSwTqW
G3Bz6eQnWJT0YurLHGjn0TiCNt5QSOTlgEoIxloIGcUwL5XxaNCZBvum282hAm4XVt18ly7ZWHAq
xZgVWOomqYXxEibl00SROnV+qE7kxn2uMCit7CSDadOSjb7M+kiShph/7tdfNe0vv0oggUYtDDfx
SHtNQN9W7NZldUGgCaRusAJcvW1PMFN868yEKwbXh6WPjKwNbuxuwbtq96S29DiowXo/CP3668C1
6yChjEu/lJDmmjm5cNO0ZDjzoLIs9Tp35ez5H1YcVcvuMUrXz1cql8SisPMvyOyiiGAx3WMKU/X2
b/322FRq4cA0muE/6qmfA3x9/xRoJvJy8K/j3nFOZCjhZUdTz4Hy8iaKhOff9EUJnbeHglaesBjW
9Ld4e/3mYm/oJASu9HQlTiGpDsgFv/eRIMdzIJiilTyAQc4cqTUQ+/4qyUHp3zUN1dYdi64WNUyx
92mrEUWCK9Paqlp71JzbDf+1qe8xxC84wDMk5SuiTZc848Fe1usYFUp0lAclJ6YjI+F7T4btkLxl
NRLXq3zqj/uHVUuaalPU5mCadttqwtdEmKAdAbrCM599MMuC9dQqatl4Pgt/0IVvbfTrvu9+27ff
D66XFtlboO8GcZGOwRgKgXS3kvky0UlAiAsbMdrH7Wlul4WC4n7jYL4pY0hLZaEOdW0KSD12yGCi
qkUShTNqv1scnUu/9/yZDnGgp7J34c/CtXmk/vWlJprix8Bg2vYfRNX915bAZkYzIpDoU50o3SeO
sbBk9fCjGfp3M8Rpk1l4YkiqnOAIBclElP8eVBuMj+KNzo0F92M9ijgvCRklfplPFIMhBrV8w/en
SSwD63v0alySbb2LnrMv9gH83TjG8rpWK7geqLyUW5aDGEkx3hoBSSzdm7q2DVUCdvu8gulPSHCq
GlFikkh8gQ8KMNoGbaOkz9t/7Lk8ci5XpKg+5UewbObZpn+EJ/IbwIr4wfNqG/RQV1gK5zBllyX5
/G97FDwNZWaiwhL+rFcmdsq2N/Hnp5RwndQm0abDzh6u2ZSapyfMWHzdFR9dE+ZBmF7Vjzz2lArR
9B3IMGTO4nlaMS/MAMaqtPAXEV0yviCWbgCEniyMWmqV4YuFOBUW3V9x4Ut7gTXaOJgMvGGj+aSE
C90cfH39equNf8WyyTWZvza+MyfifiLMtkkGi+gt+JhlP4faIl7px0s1Alj2zAEmP4bq0haD3QAw
WTeXRyPdgNPOULPBTMmU/dwqJSuPix2ylJCfmtRMDouHj1hi95FJ90XIIC+s4bbakIGVQ3CTucwc
yapQw20yJQlbKERE3RwDZOAIYOOjLqKcg+4mvlRIaxogFop3tCiRiw96mkjqE/YG7hN/YqoyZC82
hmnt9gbge14PJ378F13WjKOauErPyv0rvFJQAmfbBzJ3mIzLm/H9TZSCo/iEWqWloukQGyKseMb4
1zLeQ7VPc2oG8j/K7Jpfvkh1za8MINssDFOdZT9wjwoEwOSh/XD4gGbyJCBtScDCjmf0STIiz4ml
bhSkm//zMRXOcxPxqw24OxWhHAr15NDYZKNkzbeSpDPSZsU10IvHT0JbFLsn/n97/ALvqJLMOldM
ev8ZKhBsK2Xd0bWGzWAAo0csorcz6bBR0XiQSbGj4L4kIiOCNGIzOio6SnMyD2i6NCVhn0Pz/DLb
jXWyV0Y8/ESzYxpu9foGZdSHgZC2pyFVQ1Hvu1sSWl/BcXKDxg7y8KDAwR6Qx0pSqQ1HzNGtoNQU
nxqfF7PiWrh+qc4NkI2ZtR2HU45VhClLA6GeLYYETFkLXEaM8JN2+iqb1B/6ecjjnNGriWxvzmcX
4rNJqgf8Zj0OLcDm6rz5M07u+/Mo+52CsxCGS4FJEwZvtFP6lN1EWFwgSK6YQ47+2bINOtIQ1SM9
qxyfzGvJt0xSldmfOJUJy5Hh5mwca5NKmxjVOIn2LyrCjeNvyvxBy6ZOwTFFu0lHmbyasQjv0VfV
neOWVizNHYTXCHYtQHH82Qy5l2hwhjyfMvNFebmz/QoFat1yHy8AtiBoKGSNyJig09Z6u5Ry1oDC
fA5mWimzfmxpqj+rSJ4YNUmOIF24GNRtXPgubYghvFqTBleBPSOPv7bFf1gCK2KPtymJzVIMtZTl
3U5Fmwi2/Gw3dP6IZtksVVnLgYuvGtVgU1tul5339dZ7NW47k7gkGNutvcA7KxcrWp7LgGBPm5X5
tUPPaZsUJTovz8THpIskbxBQutoAai12JE+YzauzXHNXS6D80uqJQGr5MaqH0WreKqjpWPiUgs4L
TiDX23Gm3FMlhcttwh4oOdPBv6sep/a4McLfuFNegL9DU79Ar2czX8P1GCeeRY8nneR9Uo4SQIwt
mDtBN46s/7g9oAZEU6r/I+Ksu+LHfw4DHF5xaJAtKCCgnOf7phN8vC2jluQDOAyvjCqRzQXDE/UR
eOwUrzitHrLr+qlJWxbkoFlkhF6VMjI/bvQVm+2sazwOAgEfwmYbv/icmx23IpIcYIx1m/fHecJN
7f8iaREy9GaXVnX7VvuJ2s510Iipg4XVx0fKDrz1Wf1PL4evV/NfiWCVx1I8GfFJ34pGe2pAJj7+
KAbgXqH1U7wZpMq2XxzAUNuMVh4gnZFI58DBH5Ddghvxd7wwsL5dZXvxvGdpEdOWSpl7I97Lo1fB
62tMZsuKlqUc9Y2gHPkzM2Y905zxcCIlc+XzhLp5Jx9ETPdY1KYG1flIYgUtoJVoCAMxZcGF6kq3
oEmTv1Pdc30Pno1aJwo7ku0itAqBpQkNRjrSru9WL9Pbgz9qQTDizHHL9WDtliZMvlrb3DQ/oTcM
BctsVPjtCHV1hjk+R1UBaZDawSdvGU54QCg6PSbhp/NgaV7hRY6n+Aq4XG+NTPnvME9ZAS2WMjF5
QRIPhUORRUwKRyeFY9m08Y7QhBrtAUdwag97Hr8ctrtB0z1ivHSjLMgwGCRxxPDkEhgH6bNT4T6R
KukphDkP2PJem0kIXlCIeNHcGTroqjWBFHkBkmV60UW5VtCmp4EovKElYghNwLSPrv7lb3ZHhUdZ
wBJQ4W4SkuYWTKeVqXwgBge2HQlVHTTMWDjdoxmoqXOV/CBJvUBmXh7vhTbRqDBZz4bOemrajql/
G7mc9bIC7cJfEqhFHYvt9kJzM2ZaThBaQ+aJfV3tRr0qFep7Qd2w2tb5dVFrl2sJjvP82v0zJfsK
pUnSpIkik22EuL2me7iCKNmxiEdy7fCekWCxTZGV4P0mjqmf8rZIVVclhPY8frIbDtZfkUfjWAb/
d3DIDSttV1Ra1C6oLKA6t1zumhCYtb4CiBDePyQDsASlxTBpsEFBCC0aJCgWIhrZSROvUMRcMxtx
8stSsFVQ1N7b3LdTM+l1IQNCfdUeYFjyFRg1ua83gc7mTI2OQ2SmMdIrMpEDY9nQkoS2aXKqKV/4
kKozs0s/btHisrwxbKDHPL7PViZyKojLL5/hNYF8dWfdG28pbt1IyRzePjWlekCDs5YU+9YNrMgr
urtm9K0pvt0Na3kb/92Je6IYXvKSP0yueXqH8fCuqhAcQH4llvnkqpPwUgTo7i1EsXonVm1PUJwy
wshqznd4EP+PU2SoRYHwZNhPu4IT5QK1y9AIYkgXkB8BlVOb3Scs3Bbxj8ll121k3uSPYrz0UnvY
dpx8IRR3ePhl28SbRk2AX0LvNjcP7yznPx8PdDTGXmdbX7FxJxCc+gFJXiwLWBp0R+lgaldJDrL3
I1ERIShKONwZoCPQIeN+YS3DeyZThXTF8iFly4fn+k8cT6E27P9jh+Uw5oR4WUB1+Xuk9Ac37LC3
BFKZ/AJ7YO2C2BigUxiYnGq3E91NImqM/Az2wgVMIL+MgTxG8bnxjGqtjawPIDqR7fI6kLmDknFN
RfT9bttsvw2UKpZLtWytHz5noe48iq38RBkx63P17YsD5OEYMmA4EZBYB7mH1S7D5L9QmC5Fy7FD
KeGQtS2W62oXN5XM86E4rHH1bz+kxMqnsB5Ab4pRDtM2G9jdnxkf9PQwNTHxDGxW+3znvSrCQVSo
dY1mSzBeeKgBdgdaPU222aYtE+iMzHP9hHqpChe1jw0lpZwnK5IN69i+M9by8B69PR9u360eAyuv
T0IHMf/VtGS5JpNmBZWmQhHZSxqwTupPN2+/1n1rIZyDgSt1aHcJrUIaONm6llUdHPPyuyKH0R1a
BVx78FQtiyC8Obrs2BHnQJFEnAgAj9bdnmVVnET4cY8hQdY5vvCmJzTX7LLyAh5vcO5fEBwtQ88F
Am0bzo8JuC+5IlptHZjdr6AeuxBuCPOqspaTcExNccUM35CwNOroR9s3oLefvCqKR3Y0ZqaZOBHa
qT/ZLZ7PCnybaSXn/OpfEZeZ6YLPX+p5/Uqmc+KhV2SyOXo61AUslAl0rJzoersz0VYwQUntSNAj
E8prShU9iEzvGWd6362m8NkkvaQI8sq5aGTDYcVnfeZFK9OfZu4ulyD9J4TZnQfnFN+L1C2/yHJF
3p6M4cjrY9u9cZ1ZlxJ0QM28Bmp0QPpG/MZ4jEOQl9XuGvjKVJW5WYIVPXHUu4OkxSAe+M2nMPEi
dLjVLugs2EuCfZe9w1ccl3HoDyKYLIe2DsANOEnHDXfPrPy8BHnU7xza0bhpHaixQNnMOuu5UoEx
E0rN0TQoxHaegi7ukYFBI8UnrTf0lfv6ISYZjZAcp8wuz65ToFLrRLgKzBQsOiICOHpCQoppT7as
XxrS+XMphJosN9DKOhK0oaKHkE6z3ydRuwE7eqyWkbKmWgzPFlvfUjBv6Am52TV7kRkzDbF67YH0
wcjJNksA55Vv342wU56PpeO6Y8zy6c5HDQlMn9E5WEu3mKW+tIsPBlx3ix2+Lm/L9aHvU0NOpq8z
PQczOm/BgeG0di/ZUjMvg9o1H4lu1SySo3+5Fhv14J9VuOPPYbVX+fyHQFu5+ZuLK9ULHE0T5rxh
SO3JzoulrqOKc8nHBnFYgWtA1kNzGKMu3fCK6sst+5jfSmKW96aYY5hzhljMTQDFS0yDY1EuQWlg
0QMt8BuhwIofNDr4hQKCtyTmr5WHL330UaNXConukijhMnUXWPSSwPGoEWC+qPyE8WnkczLgJwhY
/WYPCS1/t4j9DyNVA8fzdyDzfy9hnGmeJSV2YAxj603ImqorH/Fc9oAoFgQQTM+eQJaxy0BRcIMZ
bFJkXoAR4LoWd59LhuUqmjjEfVTgvAFBi3nwhCshZScxTm+yifYA97yf8J5H8LVq+u+zwQtKY1vw
hWvQRpoQZLrKLfgm149k/HeL2KfO6v3L+lV2EGahNOXlNiKrpL23v6R844NGaTkP0lWQ+SuguffQ
UZ7KZnFflcYrXq5MZG9P6jJfUUR9ibvupaZUqa3SFT32elzKslKbWguu8OY2xnhyS+/seOHwsalL
dbTuajwkzkmmPRmflJOwaV1c6CO4fFXHmKVDE6TTp0gzxyL/zoUgR4gFtBRsm2eQQyA1r+ZEIHva
6IcBYpG6LV7wnO3K7jdtWci/MaNfAqoWs+MmfVAVobyT15MIsaXHK2ZWn3aUsJOnA2oVzGzmlmgg
LcrY35KLu3N5jphlQJjw4ldN67xC0nuijt/iLyJVpamGhYFX9VPDTOqsoeDr9HTeOQQ13SDAlHnl
Vluu2927bbO5BMTAV2TVjDSXjZRAfl9JN6/GpbKPgCq58fy0iApnGjN4gML30GFVuat3NJ9jhWQd
8cbRiuep+3pTKcmjUFetuL7RgrkqH3TxrSupAA/kVIxdY2SZ/E7BQjeDDHxljVASgpLLKvdRP7Bv
VIzcmlw0Q/HGLZ0Daf4uuO1RiyY8NSnpRxUygqZipO6IgHMc7CIH8aDH23i/auZAlasSgTNxrg/M
E5oDZwIXtzM3q2BIQ27hrUmtOWyZJF5LRbXDxLtOovlxEvQPMUMn7y7bRCAhLnq765UNh9nBOTzz
buk83Rf1pGN66OuH1YpJfAaHUYQIhYJJvPH5czjRoyRDeK5RACbQiD7P9Hoy3QO+wTmg4SgXqCR3
4oDXvrUk020agVDInpj9BXus/D98JbVS6bPnHSugk7l8DnHpY9HxUp6cehWPFpB18Ri/SeAMq4VS
uX0ADuoDLJ/h5Vb4LpLHQidAq2iavKe3G2PnA+SJi4mg23zdX5so+443AV+g2B849FDro14euX89
vQs4OxO4AR4F8fVESV/nnYGgI3gxzIlSzOz6XEUJyiKGcQJ/78lG9/+zTkPn3CzAfyg5IWNzQZlG
45X1lewqf40cOJSWZYkyb/NNY9OplcbxZJ7BJPcKbEX1INaJz+nP31hiBHdjIvDgRObBCILu2HaA
PyDKZKAY43Z65mj9+WHoWu+ucqkwzzdRX+GIGwKovCqtu1Q5o7mu/3OQLlMyG91QoCIocpiKEOiw
y3VETTC9tbu/biORGqAGYOqP73ZSQq51dNfxZqqwGDndalfEwUcGkEAdRrtQ6ZtgNfemlpGvU7Dd
v58nJcbcSNDzoj0znOm51fAhp3igrMTSDMf13W17GXw+9nlDPk382aw8gehunljGtCZB5qwXqo8a
dBdqDYXlV2TgIyCoM92ScgKL86XSiSpr6AYZajuuSLF9vDjyt8Aubrwlca7CSAvT13qqGKf36PVV
CkeFxskePNQtcrMMDgkolDdim2lcEtokcC6BX0EmV1IMfZ30vx2pIQMGqILEEO8TgSC6jysPbfN5
l/ibWUYhkokolkeXMjyaCJLLSUmKKdHjP3E9Jb0zPZhukhDiqwNwdhmYMw+f3qa5BWgza20uv9uI
4cUhikMHgisgtRzi3D+IreZXuojWAQmdGruJ/mzBkfZ0m5I+u56YtyChjtFQ10+z2LpTpv14vmGI
DmVx40Cy9YWBUMSLx6xaFoYLuKdYtfNyQKjJiYJ9urLHf4doZgbb27POgc9v3v/KAioToB6bNw+7
bR0zWTMYaz//af5sn39sJo5Ffmuvn2b3Mhf1WAXlaW/3/xBXkZS4c+A0q+MgBV50XuqiazDOQPLz
yA1j3BoFHw0MIHw2q36EieGUx6PVqN0cHlHleS5rJYnuqq7s0R8Sa9Vae1vFUrx6yf7FK/9yal6W
cisiguFEqGtL44Ig4Frk8GkN3OGP6mqih++16Rqfh7XtlhoUq9ycPTf5ZRcdC2RG4hjq8LT78lX4
E+BeTSG5Nc/ahssgx3eCiPV8iPDY7FdX2ky2BW6EnpiIjBlNwqWrzfQGpyEZcyCOtcMGEzL0qxje
qsyGAhx9gGKBcI6rixRhs4Eh9HGp1ZdhsX02XjJ0zUFZxgSAfxbOi65mgRHBHmnqQkIn5QB2/n8i
Af5z/FGeXELA4HZsmq3FSMTo5sjM0iOaU9tAYwiixq7hLtPzFWaFqUXKcEQzf7vpa/KvTPezDkZY
uy54ba6ZDyGAYZtrSnmu5ISnLiJqFQU9lcWARYMfH+25OnjWoHDH3u6r34wvdgWvVt1o9hyOQqLn
7k0ialWDk1M7jMn19kYLE/uYAMD46H3Q7DS5V0dpGi3rGXpPhfvwcHSQvx3FGJdjjRAhqwsiN76E
c7McS63hkmUPBI8DyagtAaO86NZtu3R/dqt/+ogbJwrzQZXzKv5Efu87gzJnlDn6Nb9sNhIA4HNL
ZuheKUkFZknnVr9IwFrskFBAen79Llvg0m+2yqvz53xmLQcAQ6pYcnDNTwS4884uVSXP+fAQGZ8/
pmVevdlk005yY6lqjdUH5D5EmKuNa2WljzTnjZSG0WyHoPMzap9DLUclglvZLEESDHrufdEmsx5v
YIRMGFoWFRpLSl/5oTjA1pJBMiliRl/4UYcSJpBE52LhxInzowbxJwzkDascOut9s/QT/LVN/ebt
w8sQymL4KxhZAIESA4tJLri1klZkx2sY/4kV9mkJofuRPG2sqGyTsa+DRy5h3yr7H3rbeuuOxHst
7X397GKFosVb7S6mgfduyuD2MsL9E+QBYL3iy4Fj0yO0yZtwcwIJFVKW0F7vquWq30yPKiDd8e9u
zKHwyzCd84gC4O2CIfqVdLmTKO+JxfSoFuwc2EsP9FETVy60RKKKmoFWS0vN4n1+YyGTW5uutVtJ
xQJ7P5weeDNrUcaWbuC4IxYqTi/BmvOZWeA4ZrqL5Z5tCw6IZYHhCJkTDWvQEY3HoL6tf3LU8hxA
q4+LO21zC/sraE543jZboA/DJbYTVM1dNP3iwr9Bf7m8rdRcESRM3WQS8acCmmalIEMuAyBIAepY
F2zZTaUxwOd5BCgPQbeBemcuXwW1OGS9aon4lCLeND4+t5xm0xLZ88ZFCmYpAxGzrz/QJpAAzoeC
GnuBLA9CgDwHoBk+/zVVsj9fkagbsCJAbfBFDlOu+8KRQuQKXcLICriLL5zB+AdWOEnPEayZfovy
WhfrA0WY+QP2EcTYa2A1tOmDIGtOiICVerm3PeRyBLNR2iYkKVeteNZkSG5soSYRdaZ6EFLeXyMY
H5xefFma2ti8J5mG/UyskY9htkdK/hsqZ+dGvztb5VgUFaoNH5zPJESVFLnwrhsfEQ8Hya89VudC
XOLbPOdUw79+ag4Vk4odgZ08KWIwnRdYyduFyCGkBjw0gq3UJOSRDH0dBX+yWf2TyWFV4eDB5Lzi
G2I9gIHfRBnJT12wgbGhmMoltatOJ92ISLwxSW/EtralFm8GkzQARHwPXBm/EHzvKZqRl3uCLbRk
x1usBMgSB2cQu9fJc1+cIewXOq+x82+aHw8VFaWzwaH6FYdS53Hk7oJyrRrztHL2/8h35Vio8/Fx
CJ3DFU2IizOUcVwAUnAjUXvMLZZOjdDWL33xtwBu1Gq5chM/mTfjO3+W9cD55G9AY9aPgejN4ptu
YbEYac0yKUzjZxZR0D/Xt1UI1asBWttgwDk7J9UdAX21AZRvOxT3Ubfk5ue9OZB/Yx7a0uFLQV8t
k8UgnbGoTfNoHo6p3awp5ZVsdc9HkB3lrx31YRsUiW0nfGWtPqAG1+pYCkOkezGsz9txmbucsZWC
V5R2d8145f6eBcV/AcX07Yq5vr8yZvo9ArsSv7Abfi+MKJTLq8CMFRH46m1JeJv+9rqLKS9sXKfH
JZSJvusqfCFafLjBLVVvbBxMG/wgvBe4HcCI4cNFWPdg264RD/ynVzFej5nSBAzOfB7FlQZeoE/i
45/uXaLBnW1S48HDLR5xfOmZyxJ28xzD6RBHtwB4/f4Xx3lZhpl6yEMsBkgDE/5hsI2L5D3k0lr5
Lzx86qSt4dbzuwcurgwbmllMh13AMr/hjR2GUrb0oWlZsnCC5HBH9WkkGm6NYv0+p1NuSg89OLaB
+Sfj+Qw35oMKU38OD3my7B+KtY36MSjSk56JcUW+QkXAKwQw3uT4EERMUdBXDR3SBxhG50971evV
DGEEbSkS5m9hSUwq9O6eNEwWYurymt8H/8j9Og32RGKICoSFTThG739XwRe2hMIS5d115HER28pf
TIPa335Yd4R4qxfb1S6s3wH34qO2CxH7QZ+lj3gYCbwYXbNE7BhnWCj9ITm5TJy+5KG8jv2lTEiv
KfjNdK5MCLZ/x9EguzDOqYueil0UGF6oleZ0N88f3GMC/VgSrGKRYhIZEZOKKVXkHsUyvKOt24Vh
uzCcA0xy2MkvxHXyHugTxikLOlOtEmjEbMt0bY5v+2344WcIckj7MURt3R+m2vcZRftFq8R+gVPl
JYM8VwFK2W2d5Vt1BqWsJuGOd3Q7quj9C59GenF5RWeQ7pkDNOQcQ4nvwLG2O/e6uSpEnlbHbRsg
A7KtNIqWMAPS+uukaiMkBeky90upH2UW233mzY0si2WQ3qwUkNgaey/BJdBzGqFO6MVA+q1aenDo
Dnsf1DwRCs6YuX0HLgGdh3SA4T2yp2GBgzVDD3z9G/7ne/MKGZWuhrY+L23a2VFWRWs57xcoUk9T
39tTJx9romBu/a81GYJio6y2he7MZK8IHEO9+9AbwWEkxbUALwaeGchuEIo/lbzk2k2+VuMvrIEC
QgBKNYn/bNVonaZipNmV9TDN3F3BSijDoEYFsCQu1MjEvup0SsOlirSCtzGX54LjouQSU4sP1ZE7
8xTSFZjMDqLl1ZADpGuALXfdKbiQXrknB8t2KHhtrYkBk/5kBaJvSvsVyVnXWg7E2ndPJcS+DLIG
BaHPiHrP1wElR1I63TfG8XIP3KSthWNatftGmDxmrTCA5YfeYCqWk1kUayEahER3QD4Ok7/dK7yO
wTVwC61evvrMbq2uVjeVAKK5Q31g80/DFuk0QCHYoATdYUdr3jn01ju8C2R916Ir5/Q1mwnjo88P
LG5iidLoIag72EABIJszzlVAQ66DVX+FYBXYEqBAwAlUZkGfYUA5Vf/qGE1kd6fEloMMP+4tWrrC
J2EuumSP2uETGA0C9bSJfSVA7pdSaDVyrySVbvnXToCI2SeyrF8QkOTy8zLL+WYsxe8gz1dmSl2n
iaQ7hy9JQcF7k0Ow4gd2nmE8T2YOIh7qHrMSmG2bDsduk4Y3dk93nXxnO9p03CDuPAztDb0+R7lj
pMn7cXOK6df5KMej0vCtbeuUi2Zkbz6Y9MmfAKcr17CQmH1xM+UHdE8UQ8UpiOALvOxw/aAfpfIC
7CxB+YpMrcRU0P+/BY4lRGRjbMmk7vw/v8VaA5V9KQT0L9QZXNEbD9RhDprpBjOIZShYdWRmLrVP
0/OzmSyOmicNMnr+LvQsIlcIgSLLUxkGRdUUn9a65FXvi0cr2OMbydlA8pZYfgNW5Sn/maX2jS7s
BWKGIWKiqm6iNjr8ZQIINEyvjvIW/nSwPJqVfyyvqLfiHhRZ+oa0RtuaiICBMg+88i7Hx7zAI6cp
2QrwHlvt+zYrUklJrG+kBu0cUKcCgonmVhiVce7J20/OQ8GwCR5Aba4veOOVnOsNUIC97UOjRzYS
fqZj3m9Anw+Gy3tfTVXWmIaBFXU5OWaX8PDq+dUo33VKgviCNsqlILJvlFxXBo1hoOf4Eg6F+j6v
ZRpvfrQCOQjlg6sl/JfBEVjpEgiD7IW6qPbK+Fgl5DWCl55NZYWnpoFRznMrRCKZvTvFdinhhaSJ
pqMYL/KFqXKW3PcjJfqAu3dR3hTMfjp5XAQff0/qP5SQLtYhxD01WsNhBTauPuZFqrp4UA6fPWOz
x24oK+beCTiwI0gMbHMg88G79IISddBq1fxJyvyhoId6y3ECCrRsK/vtC1WJf3UXGXj/X5WxSvIk
ediWkz41ddn3LeuXFLpZSdb0Qni8BHfPFPTEYQA6PJ14xzohSTThHui9d9ryAUUUY0LUYhsF7zH1
pIXTiNE/LKc36VuLvNXmh7+cFh2LWuECuoAu5gU22M3zlWeB7gme32UzHBjmOpLYf/14I7DzCUIA
WdqF2SMzaDiEFCEJZswN+U1JVTCwKeinE0717IxJ8eDu9LkKiMOhc5njqN+gAP8ZpHpteNroZbcU
9tLEbF+g9hkSfV9zv0V9OcSdZS23hUtP0Zr0dAAF5rIRAiRGaTtJUfL1dWPGEkAc6Yf5EMc66Fji
NtMj0PPjS7rmg4xMMdImwLO5jkGpCTVUuddD/ceSuVJTTs1x/Rrx5a7S+IHDr+o4JNe6iViUL4IZ
uyy2tSGRgvEfwEvcgPZu2tJIVePs0Llz5dwc+jCp6dzVgwvN/jfi5kjIZvr6biVXyvzZz/w4HLRc
zI0yiPMD5l+/TGfHvLaR2G7vXc/Sd0rPmtrAlLl8fMUZmjSlNurElaJR7BtI7GylPOvhNi9crWwx
PPPAsFWeY/9xn+b/zrbpDy7HwObG0NB866CpnP2R6qGN7wHmngOuubSAuDPogfgtPRetxsUgEPB9
2izyhMI6DLXlsPGCjlgsdHm7rfZcq4pTF2dBnzqTgOb8kOmkIkAGHSP09CDS2L0E2il8OejsXabD
Sw+qm8Frn7Jj2Yedo81kM5ir9Y/JIY6wa6/MVibZ+tQ6qMVvZ0wW2ngrVh5IQK/BZEDQd2iMa4hC
1516Ayusrd8bA3MEM0/PBzFiLBBVJLqBvaFBc8/LhGZjl3KhN4m0pS/si3ScqvgHbf8KwOuKzK3E
3XT1c1dgO8K7DeX3zGKuFAz1rATTOjUmjAEJAw5RUvhPYRjpYudbEahnJJS94aJhGXcMoRBtP/iJ
RgVHqrtuX/DQsalcsHXabe2DjZewDfwXUF64KgOrcIlTywXGqpBL14aHbsW34BHXh3qopPEX5EDC
Ou3d62C2UHHsh4luOxD1ZnGDiincIWYP/x05rAYWa7Kec7uG+W19PgJIvXNkL0HpfUCNqQbFrQjM
W6gszO3gS9sQojMPV3+gFBd5fFezlih0sfuvBalaxOO8ifQvYZNN6YulqzJYn3Lvdw85zGVRzIsa
LJqqVHwafLbtTdFBNhVtZch57z8SvZr4M1pV6hvf8ttfrcU6MGEGr2/BJlYE3nY7qAcTSJdcVQxC
LaYPdnUG4cviRPkQlBCAdLvzKG/fgp4Erwx/jPL72B4zueUIhkFPFFfuYSEZJZUTt5LP/JOlVLKT
6lrZatNXGfZFencLYIvJN6QdsDJJKiWnkGJ2NzqCYtulvZdprfEyFqvsOBFanqZLNMeNTpuAxEfz
gOLkhaejO3pz3oQ+HTH5CRxL3MjJmMHXMxNp2zFhEGKtfn81l4EbH0ZjPNqmEdbdBfSLc+S1DI1C
iefRF3dv3Y6PQ50auR7xQMgQIoivU3rVMg53W47+iYZ6wjQuwESY5xPPAcx8tEuuJqS5POZtHF+w
FtZTh/WnvO8vdLOovKGWWVsGDY2P9aHnhzMz/rDZ6/f/mYWVv4JyNT8Pc6i30ugL8m/OpdBnPWMC
e/3xnYPn0QtoauQu7FPHV5Ik83az0bnaPdpNHoBRz/2mOY4G4z4zHAozDPzyzO/BMyLqWNK4Oi3I
uLTDH0ucNH4uzoR0pFJ95aDydbPo9yvRHoVTPG0xRqEV5L6KMgPTPoHGshPyJvdJmS9ViCjbUW+l
jf6pt8y5+2wehx/VRC9/gXvgWbLdBwQOcnFXLm3nuv2nwgsBXldXFNyLBvgyzuXAzkeKRJ4bEVj4
4KfJSI+aEFHnLO0t6aoq7tD91njXUfqFV/YCasg5xOvV9/7JUSxNev7wiJlsnjDh8SiMQFfSPrMf
j/70iiFXS5WoDaFd12zVS6fregB6FcustcytZgYyJmnJUwkQYESn4YTMRJL1ArfYCZP+5p8GEgZk
sL7riAgEeIyEyALSCuMv87ZQUaOjD3/J+eE2qqpId5BEJCb7I5Nz97l/+E7SPn77xrMvJJHkkhFs
ZTMt0hPGBLSKHPHOn6UbYSlHmKUD2A/RRFhzpliB4aat3jtM+ZgSTiu49HfaFt/1M0BYrACpL+oB
3u+rdjJ8mAZfRjJqY/ack9QShoK18JDPR9XKGaz7ub0TfNwztFqhsfKzuJQiyhvpSMh5atUEMhMY
6XaPFkg+k6bKvYcrV/ORNB4R3Tn7z0G9p4SaBSKO1Aad6wh3WLhAfJ+lQGLjkGJIkfBE0zYaK7VH
q29x+P47VkzLoZgf8FN0M/NRgVSYrU+8eWmKCHoECdhsawq1f+Fq0SBXqDnQouU6tPoXSKtZ2aaw
yyWxggFFGFYJlLUrCGScvebnU0kaqIGm+8xvETCISevoo41Isy/fjXF/kKDZNcGdev5GX85eGDyM
4It32IOyZh1aAq6DSdZKZ86nMJox2M9BuSqFbW6CD7jX6c7tTP41YClk1v1B4fBS4nRJDEqClPe2
0c2gswxKbg2JsvGdyKsEvSx1Vi0V6wQJ+omMnZYrFoGrdgAhqh3/YBzTDfpV+cdC98Jfo+i3MA1k
MrbgALUSYzjVP012mguQzSZi6FvDPiUDPS2Q3n3ZY47yhGko4iYb1fpbSiVSycgRK4CD7KkT/rjT
HufiPlwQ2oUbLHGi0s3sA3zV9tla57zsB8DolWK6Mw5S29hgleSAjA8WmLr58DCHuw284Kw1x+5t
G2qlV9BGMmu/UctJq0oOH+2B4bfcipE/XUiWHn6trd7VBlFw7Rplmpf8eBhoVZEHXsGg80g6Y4kg
pi9MRTWvJPI0aOSgAy2hnU6wX80bt9fRoDcutYUFXQhJofZ1CqqH4lmbnATjmEV2M23jxOzKdaCQ
Lw9q44ikX6AzKjYbvoycseX9qXaSXveDYPpT/yKZODkDOcXIV0mO9UVw+n2HzmrEGS4kBZFfD1dC
VLmMgzdMlXIMG3CjZ/swj5qX1x3dS/3D12SF3X3u6xqD9uWavLM6/pHaGxqdTdupw1VPndJLT3kT
Op42DcANxVdHpeobW9iB2St/KJAiHH0XZxno3WGcYfc5ytW25bgW6ygYCIxLDh9/WE+EhMho1da4
RExioHBz80zob5HLCD/nZB/PC1agLFA/lfZcxqMzx+XHi14KqUK4fUFhTBosugN8Jzz2+s2CKfTj
cGwmWzHh04XMqIyt25Ig9crf+Q1+GxU7TbxkSIM5LpIrCbPPQKWYe+JKjxW5FCnDPov9X9V1GmQL
sOPN2uxFM99Z3AeueuuCQZKeI04WbX3+lH/TQYTlxmXDWflfr8bXfFoBtRzoxlObsTlqg9XR7G+J
9r3wt/2njbMYjNH2xzULnAvxGVsWmkFV9hZl8kAqmkCYvoAPOkJpshk8e3Xtx5gNzUfxuUnlo4dQ
Q9F68K/OGWo7oUtEJ+VyT+tc64oA+b860HGyy9m2o7K5naFu/HNrKdxSmamW0dxa0rKmT6kKVubN
45pTY54EJJUPejug5fKl4AvxfvTYy2MSBVx71VnqfG1J+qG4jt4idoKnM2QxuBNHIsrwLbO+bLVv
EU34XCYUNQlHSQFrs67MZEJwQ/KwDPxZjKI2gUg6ApIj7iMurgy5vVVH240rFcv8dITifT26HLWQ
J0Op/+DGmogXlGxuJuIoEDzOVCwyhaJYXF71e/Qbnccg3sFs8T6JMVPesybXlnYlilk0dfIf1xvJ
976WMZydzazQ37zJOHPZAPw1hgveMc0hnHkaQxcLwhWslP+4zTVTbUHddD6LQhYFOoFD/Q4cHZrc
i0KvXBNvLtWsasoLXT/L1o5OUycxOLjSpFAYJ6DK8l+LOZCsmswP7endxcV7QVpTSse57rZiotqF
pUYf79Ln3d2N4qucmoii5MawrAR1qEWrzCrb2tvX1BV8NPbHyQhTD7i0KxoW7nwH+jWbMPM3d33A
bOh7qQ9SrgfS+3caxRosbeClSabE5fs2INWsGSXFPEMQjZLxc7hMRlquAD2PPbQQofwT7V19FyUO
WDiMvrUN8BcobRdmVHxelNplthvyceYE9QxGP0QwaK4jFg9WV1ueiYyykFcKSx3WO09HaKjjRzCS
uRtKRcPkEMVAUCpgZdV1YMJqUu0+W3IoI5lBXHM4njQNEFU07TmMCkxiyisWYJDDZAeBCP3IY4+B
J/SsOK8NyPbLdXn2mmT7MfBUJ7UcympJTIEXB9bscDxCS2w2sR/Zp5HWw/rNYXt8SCZCMHcN7bRA
+ZztJtMVs8HpFigtgLZ444aSYzcTKbp2jqbaXGA2k3LZ4aKzSfR8QyC49C1j6yImr5bW7L704fge
97EfHmL8/fN6EovAyfXBuKxLrDO+tV95uS4mlfibi4Y5iU4T1gyDWyrZ5GM6RAoUBUzhh8LyEwWs
Nz1xaICYpmGAh9TtrjiKq4DelgnW4wRbiz/ms/NpmJIegLWhCYNKcytC1XaBKcoCOlJYR8s76XjW
Skt8oBjB6ojPIukpjucRI2m9Zqho70KqeSYX7UAiAy+KEKoIGXi+VF5tvjtjks5DuiLentGuxyw5
2ZB6zJKV176NsvMwfkmJ1dd4xFWNpUrJFDJpzmN4Ns0WKQnFgpI3PHK6k5m55ysS5N2lbECmRKbl
bL+OpTApDjIcklm88aJCiLqLAdX4ql9DMgsane5SDkuCWzAwccC0+Vt//umQFDYicWlIfyCFfZBj
Nvyc/y8RNkWYgaaXE2FvrzHv1fRD+QrrHNgkXfx/5CqDVSjHEM12jAozIotKbcuenOXe3mh4aI0A
Eo/xvUdurh0iQSZEGTWv4+oefuemgE9L/3KqFfSM+y/s0KP4gafMlH7Bv6zCCChyTXaGhIDU/g3I
mj5ZwvIX7+BtVFs48jx9KTrYmq4tPcrLjUVEeiHzgnDvyMz4B0mVPUOmauJXIID3w4jjXI4bcFPX
POD03R6tOhYKLED1POABCho2WjQif9EpBNPn1ClqK8q4J34yCa/iQHkXuRbSYooRWQgQJiqXNHmN
8cvkwIAsvbmh20yiwD2TwPDIn8IwzpaUFlnfPir2JTNx0O1pOwYWbh9HES97IDe7OLD96hfAfOi/
dBBmYcuBD6whh8XsMBAOG0z/sVMU65dzXs9+qTCERYTTDxDltS/tQ4O7koGQFVdsI2faBEiDKIWI
gIq7SYiDwtxLLV4Qu8QgcmRRe9OMj3748lcSj91QTA/2Y0HW9z6+E/O99AxncBNhNQM8E21g/6XO
Qwu8peWnM1enQ37sb7uZ0U14Qd87gD7rQwTDdqybwdYmTOnJqcW0/R0cXmqrbw82zzq1lHT66s7x
Kc4kZcNWauuB/dYef4PvxvmAvskDpkI+9Kw3nKQ6hIJVnIADMra2MOZWDUTNtIiWKrX7nMRFHW1z
R9HfgHMzW0x1mMKQ3SaACTs8eQUu4IsiYWZo9cykRnmNKY00tRl1qeKxG+PmFUeqRM/wq2QeXkz4
GGVNGb3UrVesekpwEA1blBZRf1s7ABYrDj0NgzqUlzG6EY4TqgqdJQflseIyNjRHogzKTNm905fN
rrko2cHjIGNQMeJQrRclkkQXhI078uBB74fspR8hXfTvegajyKVSfywsMUtCos5H6OFgWs2CLR9H
KenUAo5TYhGpeeN92+0oT+26FUfU9uG4yrXKGbNqw7vthIpopSfBFyzSdMOMlnN8XWtrAjK2r9pC
8cGCqdvQF2J17MJ8LTEs9vCV7gbIK7ixe+SNDPXKPiHudhnVD1BkGtQ4ZrHh1otT6NOk/r3eoWkP
3ygaZklfzGf2eA6rL9m1ZLl+nxLrfjqludDaioQYq90Qudnj0tn00DX4YJdD8+Ky2ZpKPxu5wUyM
KGQfXNqNbXsWZP6XLkLUAp9eVq+At9GlEIxQy//SdyS+FhH/1lNN6btd9qPIDkL7AI4qqGYIbXwQ
ctSo33+YxBVr/jL4MXwWsSSGi1gzscOK8pYpcxHO10A3En7x6E0cUPibFqlAeYUdYQDCU6lQ/Jm7
l8dv9xynLWHDQlQpy2GMaJ6SkCNgaDMVYBFCltoP/OkvathPfDtST59lU2s3cdgOd6Hg+74UluCs
Zr14/KfhZZj5hF7maXkP/nq9ZM1Mu1oWmclQUo6r8SZTUHsCgnq29dT6D8K0fbY9tlNSrn9O4hHx
rcFRvRUSOU3cp0bFsOOu97iZj2UThKD2haFmQO7CIPZzLb2Ei9/ZRF3jyyh5Pq8wWaHfKs+WM3ue
V0AXEsIaPGghjLYtUkpUFu70+Xr9vRFAJASa0kJQCGKFUqUhQ8tJ83Xs0BAv7Zmhb9LLh3eDR6b2
y+3HvlWfvYL9yXed8m8mQId7P4tv11A8Ts/+5yrE5xTUpmHnw1B6g5yReVX8eqvexXTsMMdEcZRk
zpgpXGH4zUcrnvitz6z+R24w1zGFLCsB4XQaGf+C9qJg2qCuolzXH9cINzeSDsO5QmYvkis/mfoy
5uBp3ATOCbnCQMKmT9JbUYljfLxPu8xGEKM1m9TG3PPOGGSfl9xbpcoKGJ69EddJg5n7ohuN+6FT
onwmwJ5bXV1bCvPQT78FiDWUudM7m66VhG4FtNtDi5JuoI7xUuh7loxVKKil5mxW4AjzqHTJex1l
ECJ9sCCouZVMPah8hhWa8R1y/c8X5v1lVGnzgCNb91iprMbBTkcDkQTxtydgSJnsf973CpCmtFpB
Ewe5b2V3pIETo+Ok+X7o7xFQsVvlsBhglQ89Fw34ek36mkOYKJFMGZsV0dgOS7t5NA/Vv1oKbcl8
FBRQ13FsX4AvK2VLttEvcQJws8pw6dnK01LCZvdysuF1nxMuDwXc2EjUhO6rFj0qb23mR4pXqeS0
9QWNeiYGcbbHOZoO9nQV7mCfMmzV7sgWd4OqJY9H+cklv3xqjwbfP0ZJRKcwn7RSwRTiEJbtDOTp
XQgjU9eJyPcmQMtMwNfo7xquhqfnyAm1BfSyE2ZB681PZCcs7cgh69eG/6yyhjRErnm3jUMKMX1o
hBQ8WsK5vqocbzjDnQaadAEbj4LZYjp6Ne4sHHl/F4esBXnwiToZ/IWsjAQpNKPPywNL+tGgx3vf
QTs37wlMF+o6h9zt2VigHSV1cZJL7vKJk8pJp/kmeknr4wOHGeSex0tIqREeWIg5UFWTi+ilEZiC
v9jRlqwbBz2wigfefj6pau1Y2fcshMCTiQWRUAkoJz9OG2WLUWTQhtEgtzJgZFw7NT9czagi8YsC
bmVtM+3de+m63ayeFSdOZlAGv18QKBWN/OpN9T0vQjPqwyBU3D2qPDNCaEtTtuZUMQtplVjvNToH
YzwfXAqMGfpEqQoDwQIra/YyVttYDNiBHnux08rblA34/9w5FpuSjf7ub9tsC1YZJ9NFOX9gp2Rx
mItl+HLS8spQURH0LOcbHFpNVdXIq+Z7SOhL12GhNwqV5biH7AljEMMVWNI1se80yzvJ5f5vFAuo
br6lu+M4GbPBYN4QVZTaBowhZe6qDRDtJWXDQ89z35nGizVYi/hBsfz1MJFe5rITTOKEXfgGAxPx
in+ebP29MRINBgdeF0OyUcxS+Cw8pVkeHX/Sr+RL9TdqxlyIMAPCGBgdn8+au+3IecQ+g01AILXX
JMYs6IKgpHwGlAhVrA/LhlaykkvppmmNuwQLa9YoXA+jvvU3yvStvIpyDM9EQPuDEdGfMuhBxsBs
/cGdTK1/GhfkYAsM+tEkMmAEKhrIZI1rFUGiKVaJnd55pkDmPKdOcFFAqaD/91MMwdGUuHQdx9Cq
8ordQBwtgf+6S2yQ/aX6sqnKMMo8RNqaGCZPYNMHwrpP6wX2BhOYE32OO/jsrxkwRUU8FYRFIWOG
yrDb1tR+beZyKPvSyM9TyVFLfzhC+lo858hhW4PveCGbpN/wZtxOITQWzWGVU9K2+MwtBUREAMW2
gTmaXoXUC9KpT5Wboo7FyneniNyKYYLF4sbRFIE2TvY5QpfChm++dZiSd+/v1Re1kaSt5MHT/Fln
0f+C5/4Xl6TKsRQ6vgSnRcg/Ofk5637zc2/zrtwwNtNT+YRu2wkx/6EfFJdGIr9u48Z/Xh05t4Ih
WTiz/Y1MujhI80HqS+96xKRNifZzC4No7snBJawPJd/5gM97/vTrRiKw1F7EiFog+mP9fJ8TVvf/
K2VP78emijlYHJOE2nafW5TDQwTfjiHcW1Fmw0T1cZ4LjpLSAPQt8TIKSxsd5T3KmWMj1NENz2MI
7VAJxbDeCS50gl7/Kq/bKGW3frBSTiNBG1/Fg7QIjLPgjA5mfeXjI3MEeQjor9196ZZqxGV9E4ox
Ky035WlXEixjaXLMgDk8xv/RA0KljFx7IWr/5tq5qMP9ianWy/nKOkZru/K3SbVGC1c+7co9jqka
32LvR/oiT2FEPLX7N+Mgy5I2tQQA++IwxWwhuCHxqHhWJoyDYyqxVyVwMvzGWwtZGCdlnXZkIWwv
iuwO0ln32xsslldZUaokV61D+mzYbF4RVZelFyp1SIizbBvqayO4ZLcRg/FkHIJUFhyGWoNIuNd+
45FNBiFRhqPAZbbcqVC+EF/DtwrPzQqze+Pejy7ZTqwleBLSoXxQI5Ar+qQOgeT4cgFroOVERxA9
hVABG99va67bLqvnDC/GQpEaYdda/eAGfUM5g5RdtEGKcmk85Ro2mFYHanhVLnLUgpwF04qQojZT
xo69mfaW/Xae7RWhlBACWSJckJJ0dQd2LFnC/BbK4dgOQpYb9YaEam9J1/NDk/Ma6wnC/T+fREIw
VZ8rSA4jvEFsJ+JTmS4zefinIGv28rMvEVXN6H/w/PWF2KT6ysca2sq8GlQB50cJ52U2jRzbGm8X
dBPjw/W2qOrIAHExKGvbFWRZs+VruuTRVEvA9t5ygpfQVANd841VL1NZYZGIo5Ww2JmXVnT/Cwk3
FVNIn6h1b//rE54N3Ob/s5L0b3YaacbUwDDgaPBuAVF22LSZri+YySa/H4Vvf5arK23u5QWX2nhw
GRUxZHNWrVXeUkb/igtH+GO7IeOVyyMYRB9VC3EYwWt45oQ4CM0AAsW2dVqkBbi8VTUUpI4ytYPG
W6NMrQEjIedljOhW51FNuNZicM8K1e6hW9nr9sXBqnoc2S2+Q7DobNjgB6aVY1oqpH8HQ99bElk0
dFjhuV+Y4t4VbWps3t+Q0sC5lxGojoO2eJfZFV5qHZUfWx5vgYwd2aX9FXl8hbcAJl/LYfKMG5tA
rkXWU9KIaWRJAFpSD/9miuJdZWr5sU/QOn6/CBlmIlZ02Dswbf/UgstK5BBz6b9IGrutX1LGInKp
9nI7uyDIuwiGdesiskdDrA5DIEoVPbG+efE0T3PtrBCinc6xh+VOoyDfDMnQUJ/ARH15HIbI/Hx+
0ui27L4XAa4X7nxqfqh6h2IqUVTIZF7nclT7kzMc2GNKsMfXvUQCjWrrdpI+QK562ysBrJPl6O2p
m4TiAJPMm4KSwZFRHsjGRq6Lbcik4G8WQ5jOQvyR54QGMG9WG+wS6jCdFcRiTfd0uU0J+0UWVsml
miyOgCvJ6fewvlcd2HKFNONoady4Zgs9JxG98fqpybnAM2kgDltTxvaFFm2pF7nFFhupdExFVH/M
AFoR7sO0lkey9KlwR80u3NWjbxPkKnVBj27o3Otkj739TQ0utbLFINyINT0Ln2l3RHKn4CZpe69h
/gNeS5RzBa1yTc0H0c2ea9joQvzJEl23usUcy+ida0VHQGzLeUa47w8TlFkRQWg3Z/CP2sGE4/wF
fN9/1Frfi/kaEugM/aEHfwhTwg4BR6uy0ov6a7i8Gpp934isg2GJF1FM8GGygR0cjSqa8mMz8RhY
FJVykRsRT8mr4Y/U3FAU682jNs9R3roHa4Cu01BQSB9JPmR8qGrUmKcPuhXiReUC5cyVhvS4EzCA
wniJ9m5GH1YyFva7IL5TbVGu6jOdi4zoGEQFctMvVcBmnCyU8Lw+LrnOYH82Uy4oDF8SY6hbW9dC
YVzp4mT09xKNTL0coTwRv8MEV5o1PlGWxMeY2bx5rQuvLy4boX5vgBBiKSWM9+9NCHoeopLIJ3uA
19LNBHYtwtgGcCuAFrPjU6tM9v7jgSLoE7h6cKI0DWmj8rgtgHXaraXXsZmlo4305z2A/SlYk0O6
KR5Gq2g0fPrzW6oJyQDR61I+oRKHLJ74yRo7W+nESIMSkxXx66FdomIThvauK9AC6oqi+z6LK0jW
cZ4sb2vAelmWiZ+wTCirkkFq51UPMxu9BfoaYKZWoaZb0ljLWOgFxdQkcbNI1lIZMMOm3skimHy6
npsV5/ael28Oej6NibXj6Drkspmm+dWlnG9HcM7wHasY9yEU0sS4kJKBy4ZNqC/rHhwoUxLehykP
C18vR8AkfNjV5chxzlT857p4NGvCw/MdpKDuKW2NWHncekt51xa2bJ5AgJC8Pgp4ndZya5TAF6FX
7xvAKRt90CxMzH4mWPKg+Cla2OTT6UBqL6Pg6v+0GwcB6I8DTZWaNO/32TVST01tCwWZzBXDS1XW
Mc6VD1vWrwwnKaYy+t2TTT4p+U7yhMEtocPlNSho/0Wla5tD1JpSTwoUwfhtTlAwHqrcFA380DfD
jl3e7zK4NXkkSJpa2JIc2O6wtT12T8iYezJ59hkXZ9bwcBEXIYIdJrglhzjDTPlMe8yTe5zPppJy
5aMNcCv38wnbzC9SOgK/cKzXZ7trvwvtmLT1VfpcyYqRFu5orCBacIOsXh7QjXwSyxf5B+LKP6/K
uQudC0MwB1j2M3UDE+t86FvKNaI8po/aSCg4ga3KXlEYIhdvLp21d8juto9YFzpUiXYpHHx6nVde
4A+s1dbZqxQhSG+epzvP4kw5uraCi6vxt6z7HBtJnvmNHtpmkdFgwuu4JlrMcJ/6ZP/9mYiGTIoQ
4xoEXAEcShkD+2FynKni/oTTiooKRpzVDWaPNRbjcoJdg+Y/bxJn87wQfS+NOtbTD1pxTFmqxECz
RgwjmTh0BakLl0mjCbG5ax4tsXHIHG7enMicZvLMhtodFTvnTSKyNLTSUAoHN0N3VeuOvqH/N5yU
tb5eyBorwh43ISVO2DM2GszzyywsUskSY77SknUJGnq+uyVinGnXRaxoIpsBSQ5w4dvpFaEILTDq
x9Rp/YkEVDLp8yL99l0Dod2FiDZATZZ7lKV7HHdAPlvw5DJDZ9hGVcMUPEBHa8b6FeJ/V6j0Qbbs
SMg5HGBHxPvDIntmKcGh04ORNBFq2iH9Mj+B4k4WmWSwkT8bayRpwVfmPVEW5Uz3ww8oailIddkh
Z9wR1ZTMPIwz5i8fF4mXAUpAis7wbbGIqenzVtZvT9HqoqnKrWayrXcmew7RQA3QhhMNPBYtX4d8
GNoN6/x2y4YUXK773Oxpm9MbKNTRGHdsyTPwF3yKoaDwDdSdesYGwbfCRv6h55eRfyXjrJTXDHUQ
EG+sK0i6JrdBKHn98uV7pywVuby+z5Vl+Odqt0ywI45j9bkvAhrOPNa7K5tYbPHp+NpY/+X1Vkle
d4abUlwZU7kkHGHvUsxwTAFTAl2tigl1Vd0Gt2JsykvF14KyDW/lkTeIm/Mfh21Ztw+BqezZYvim
2PqX94BTmgyX4thUa01efkrU+8ncWW7rfix7Wdx+8HjEQ1O8VaGoJZ7NCgsFKkdhDwAjdw/I1mQE
d27GwSIZ/DMi29YzhLzxaKvbsjNqS/gcU3gqNHyNn9XfqMSCh+Wj5+k/5Yn4ogu+1ZnXhyaHcLP2
T4kek6hAI2EySnvX30noSfru15n6zaiMSFdcjaIy6HPVv5OFpHv+nk2ELmxgMQOaTB17A7OTFezV
wZ5obeLx4Be9EJl5c53/jM9LmGF0ryf0G6PKx/wBL0XRRgk+I63+d4hl6OWfhVexaR7nh9NftQpb
8KasV3clyvTr96M2u8nk0nhZJqC2C57aj5CcGF9Ji2xBApP7JWYaxOnDVZ4j7ZG+zZgpT+UpGBpF
OHKmelNXQJMbV1Tq49r1xBMW8P7ZG+7Pa64ll2jKyiKM0MLPSkfoEY+/YCVdMm87VbypqIbHCFHd
A2m6e4BmH32hYt0CLMbcSjxVmpCqPjKyGYgTTHxAJCSS0oxe5kudwDe+I5JQiXiCU2rdrYH29uWs
otJg7RRQzCBxHV7VraWC8aeJ81J26lFHXZolV5DcULBFRIFuTA6G6Iw54zqFT2h2LLc8ZC+7bXTA
4hLtThxYqvTkaPIesocedhs6+Dahs+V4Y0pcwtvd4NGkPeUkcQPQFqR2+0d+0gtGVHD0E/NyKOr/
Od30c7siW0zyHZ5+nAR6WiBZcNO/Ff5Td0p82ZPOaN01UtfvRIOu+6ZAvwucktFEjMW/1SLo/TC5
H5gPqRQZKDuc19gEGpQjKEfRc3nMUsHuWaqp9jRIPm25oZTvrECGkA9DebLFhMyH4D43WeXqTaG+
T7OCyaO7OCa8Dh0HRRNGwHOkpyXSwn7yiPQMhz/evSRFuaoQtJi1JtJYf95q9dCheaxVvZTd/lQp
hjtIsHo6/NIVlGdYLig1fxPpPYOs6+elj15qYqPrQIKhCxEyEPy5AsTyFejAsr8ijTpUCSjnHn2u
TXTZmcGefu2Cpf5ANUdTFhLKo5dB9swMaq3mPLR4vTre1ZNeG+u+Sx8NVKdN0tJonkkbeIucs2pV
/fqu9K201PTFeRj5cb4L0Yh8OgPkjlzBUFCko594/cwzVEpTaWs1ITsF9eunE3n6LFuThf1zge7V
qUp5uOJ4f+EmmsGlTElGk0P77ununf68ha3hj1TcTttEpCvg+kTjbjrKO/DRNp1HWmdd0cjIY9OP
yNnndYf8xGbM1cfsd305n/lThmVkxlo+R57ug5bEpZlTA7eIJMjtaaLfhEX436Xv7P5du0TXbTlF
UxEG4EEYwP1FG+C7TVPJo5Y13T1nNASivTVRdGHxIbpuWtKL4t3IhEAWk+DI64QKG5kgHmWsaDAF
NWna62v1KQTNI7rjJIIim3kpAAX6Wcehfbva2ochDOPTwzyiuiWu6H15SkUhbEHvBIYC5ncudSBQ
IqajDDV29xgFBQ1/J6UWICzwceJVgnT1tDxCvX/DoII8b+f89Ihp4/r6hHVM8PbM+tHhi1zra8D4
jzFeZi9qmtjuOlI8PqqEZj7cUlTFdKuZs0owwuccPEGkr8okyyvlpqRy+dGWNFZZLqn/jotx3/SR
AbKW9oOQ4rF6FXWoHomDZqpYRsPkfSRX2HYuN+RdJCkKOd6rztCR10vOunf6wNgCyKq8X+K4bBlc
xSXaaQ52VD+USXsEktYQ4lq5iKf3NLr5DSzTfUn47iyQIjmXf3wb20xuTOJ87ElbnOjN8rfPFDgD
WJq15SudwMaYzVIjGVIncAVnrjehGk+xEXQrVxGwBwUnVk+dszpJGkPqKcdjrygkbKxrw1LGUXME
tJq+h5gAjbsL+WqSVbHWPwoIjcLFQaC/wc/2lnBoELP7t1/HsxOpw3GXQxWpk+70zcES2XFMCz86
qmeu9Brl6AWDDXGUBZtZ8i+lOHN1sEYe+A7aWcPmUsK9L1sH+zdkyiSPiGWSNp2+ORbN6cn+aI+5
ZZ8m9UAFFvWRa7iA315WEAJOp35tLBk6N4n4nAxy2Q+B/kfJR4rI3DbcxRBW6piS3nTQKXjEiQa8
3/CHwIvsQ7MLwNdSnXfIb932r9ixfuyMHCNQOkGbrzLfiPSwDqCWGq7OUw/FOjUEOqz/LoODT94k
Fwa+qEG6UV6ZDP63Dps7FWIdtWxJxUYQB2skvkSIC2nivaUOpg9LO7cs+FUT+4b8U08blOhzCohz
K3YfxAVLdt+wOVXNec7MoaP7tQpyqhrdZABdLCGIyISOTJw0rrEq2Z/sAKQAriNj0OjUYL6YojqP
IkhfmjxmGyo/mkOKshTrlF0NOulDY44b/pnguu8lZo7islA6cWEfKiiLXq0+xxQLT0mdVhN9258C
Cr9YR5wksDCPXnCKRqha/TPyoPuAXamVqI7WnrYGX2yI2xKzlK75uaLcXWfTNSRFriBwrG3Q3GKz
3p/+BytFHZjEM30SCWBO2ddll176Iy4YXH4XVRAa7NPUWbrabONFYIpMG4aw8em8ZOETL1HQ95uW
SBoiTUv1J8djQbfHHDAkX9CgPQDoZzwXN9L+OwSjNIqw9b0VZkC6TI9AqFdeO+Cl8CYXJZ9wcQr/
QobdRgoCHwzbuesmU3dJmf5zB2JXOAnl51yKRH7uWM/1gPipC6Yw4aE6t1jjUY4pxnCpaHHkK450
+ERUG9C/CAlQF4Hi+5QJ6SWWBJ4M8qK8AUX2vGQamQDcBFVLMRzTUnmLPQhnY+2eo9JTX+evkXBT
dCxcrgnndkUuIReibg8BWnWEQpFaQ3aoddmcN+aHRH7RQf6bnprK8rd6ynn8YnBQCMwJkE1l93Gp
rYCfUgSFk//zl67PVOq6PykdX9buXALYg38XgVuvBiGOD26GO7KLCbO6lMrsEL7qv0DIPlE9w4Sc
pFQE6IffZqey1tpqZSKekpDl4C1EYWfL4ZDGTK/Qo73VDwbousoVWcp9ME/Lvc2qDyH4GpGfuBFw
l5jNf01Us5LOtuUccuveJ9jAD1hL0TX/GhZ+WoeWSxfG3J4VMpzG1DjD83qUAakSVrmf6rXKIhP7
JRdKCapfOsbYuEeYdxxWiC5TLORhAELT2q8Veeb462b2kTZgn94+usnQfLrzYg40d1LeIInrSC9k
bmRljfuj1Ti5k2p5vjzwBO1JcWGi+uD0yG6S3XptfpKbG7oK8m9rjNVm+Brwzi1vCMgFw63zVYgr
MfaRa7tUPzQnLdVVVABv7CboDmDZyUqaR2/doLctcOpGxou/9nVIyo+G4XAXtzN0Xzc87dzQNYgA
eVbOFikbZGtXyY3T4CYRjo3cMjD/jcWqI+sBBrxsT02j/yynPppI8K1uXVUzAaxwfpwoau53DgdR
QuxnTzM4MJYAJT/Ht4j0a2m4dULzIRBIrA5/HBTQPXEtwiZjAczshVqBBGpCGw8CSWwUjQn5hGOl
JwXUR8qz+1PUDFd7lfjUorkvhIk2vV4W5ErwchwdYlBcVdvXPrwQDImmFi4ZI8Jl29/o0ly6W1TE
PyFZWt4GfJwBu2+tv9eyy4zFdMXw4dBD8hcBOKxUj34iE0VIO5OiEvAErRjGHrrNEvse3HLWtaVC
m/ZYdxuJ3phm26UYyo1bStfxYeLcUFn0Ki/UNdK0Jnlc+al0jIs4c8gLr90S1aZg/2fVzYeGum4N
9zhuIjgZp/3lUJDnPAC1i0sBx61g7pXNz5guO36WnhlTTjzDnuG35JnNK6GrNR9sZLC6A/zYI1rZ
8AQr7JKBdA47hHsG4YhC2WDq89pXLzWZRehb2N5LR2nJucUA0cWwNL3pnNSa674MRVdPSNAQcH5e
1ndWL6SiNYCijaqMFbCRQRZFWtZAYR/h4JqN0tahkb8oxvLHlw6Sq5EwyS+vcKBEzoRFVvbJzfTF
lW6afrozTjZmU4u5fz+JPacPyPSrpqPHKxZJQ3RusLFDxbJjwzSszSH63MESrIQpBFLzvONEUEjp
KcJgrBTKPvAewKffUlmGFu0T2HuDAxZtJCDWjF2eqntAjb058x3UqLVkbmEVwroRIh93sQsNLk/f
PfmkiCvdl2NaZJFPDnrv7/5bX1Lulp4Th9YuhGUh9EEAJ71cr0fnvbrBTF+3zySztVemVQTWkZao
1YRa30GohQtlHv39D+W68V3umT9cpY/jak59U8ftysBoTRvvM0/5RqQoUx551juwUgZPjziESKYj
SjddK386/6k6eIGez1uq2Hzb/wdo/cihmiYEazPKT6jP4D2jMvB3co6qd72skE16GH8yl2TFwIcS
U1DgTvQhKZpDeLGbC+B1BEqEwbCQ4ZCHo4ulgySk4BaL/dBmG7v6vF1XOONpAONbcid+4oBOrBt/
tUh0DR0vaLDVNeGb/5ZbWblYgTziopmKlTdACCyMpVRjcklRLRovN28/43cmv546dbGuHEksrC9n
d5bs273mG9hYmsPm/jgU61HnS+yPSuEuAhROAyYEOh33QI1H4gE2UB5gn7HpCoB2RIiniIBqX+GB
nVI7vmqnVXt47SCA2ns+9vR1IzjtsDNJlShOt+QnghlcebxlH8xSWKH93QZUmYtyF3D99QL1YIO3
ZmHavTZKPQQdJotq5V41X/Nj89H9V2YqNeKt3Y/W9lf5kf1DpM19hMoU37P0bUmmyYtISbU1cwL8
8ClsRpOeF+HRMGkO3mro+4sxY8BAV+M6oXouqk7l2I8Y/jrUZ4oHTO/Qnprf8m390VWJ7EWd9hwx
lcVDBtmNW6RPYQRnsSQyS7ZJu6lCSuMKN19OFrE2kZLSxcv8l4ZsERmWE+X1CUk+a9IWPa/9U33B
nGUpdF+t8iF/Ze/m/DMypi7RZEEoB5rd7y325+5PKdYZDyr1bHykzN6ZG8+/oHs4u/j5EeuJXAxa
AtN031v/p7+yY9WR0OJLjIMIWw5MkDTLKbbZ+VGi4dUN7y4sNTEetk3jwz7gnU7gS9Y3e/q1jhuD
hAZ1VgYrVTQzSZzuPmILTw1pz7+5bTvm15sl69ihOu1jc2G7V9AvJ3CkpjE5y1jxUMOQivIZTvgK
rj4yxKI3LNSNCy7fwfFjFjxOWReoJiSlsCnJH1zcFtyxh8sJzCCtiS9ZiNEsfT0gWuB14IfdUGYE
7pC3OG414xkEce9Qo6FERXCUrF/LhxMYN/po1vZeblVzBnoIAYJ9QSxQh+MhVyVhXOoExhH08sSy
ZGbDt0vOil0SbRdPljFfX690qti3dMScOqJkfV9LF4ZtowJ58daRmd88cINGegg041vlRwot/H2s
GrFp9Qi9vD3PZzcosPvTW6ST6QkylEgFlt8WHgY+a51Zoai4wjiAEii+0z7SO567IIuWwKkLRqq1
R8wM4w2qifPVvhCCtBItW6/QZITPkyYlIbnK31cAksfBeXF179MfoN85QWgcWstWhLGjqeIiHuhT
nNpjPqvAUj2Gk5Nb4SmMeZRxd5vhuPlY7IwkbokJEoTX3mwzNmO6if8BXZvF1TmXQhs3U8D5AYKC
aY8V3Ek8xzAtKGxGzMEVDJhVrdjphVYpkkj8hS2eRy9ohYcWSjhmEvs2heln/RmDyj0d2GRMX4zh
l2mGvjkrSOxhR0oPKhsUb8VsCL+50fcO6JSs28IRskSLZLUFuk0MfYLveFSmOsgRejQR5VD4ehnn
7cM/d3toiH5LpH+HAGMMMlN4qFAq0lR7lv60zdlGp2nNtnoLhGKjQlou/5ubkFzuh96SRYARD6Am
T1KIYWmlSon8g8L06U4xGQclKUXYpYT2feZvgakd+55NvrSh5IbnzrQHWD018MbW5afp/vvHyXwB
QvPQJK7GlxLvycmK39xo3j6KNv6cAkVNGF/sdMgUN49hWE50C46xdqglouYPwEyqFTBQXdXhgHwV
eoWuIJUN+Ikaq0tLW01PzxUYcdh8C2+JOoE5Czu9fdUJJaGzIPdcBewpB3ngZN+O1N/OxHYonUCG
7K8QV0oWjydtrBxQSuuGOrCQzPxiXRJ8yJ8cPlc/Ts8VO3s2mpl2u1co/9GCUh6y0uPgAGwzwRm9
VnYrw6EWlWdk6c2Ynv2IXmZsOIkmEc7CE6ogJTKuVDF/gKYHRpBP9AxSrXhrlOkt27Qkh82JEm2e
7gjcMiXU+qbxSsRTU6ee+Az/b24thz3nqmSKToa7A0uMzP8JU7WwvNmzN/I31Pln2O9MA0PFolxC
Q7IBPuhlKDFmRySQF3znJQG3tY6W5axukLYdD0Ig/UYzRho7MvJfUFSijbMVtDtdoL5WyWq0svGD
T2hKKvR2gJ3zybnTRjXvqT2lNQ70BZVpUw1gdd7G/JnQjkTN9aCq3e7kVYVgz6p7/avM1LmkvIlY
aVe4CEnWklW+CiOjuOK2O92HOwMB++G4ZTIbqPhcE2iP4QdoUbqUqSw1sseXg60F3mn54B4L1rwO
KUJa2tyzYvbQ6W3uqQlUBvnB9nRIxV6oVEYSUNXMCqwX1Rz3EzhGGjXoRtO5xgftzIjfW9CBhcnP
eMyKT3Wr22qkDKE0vetAqfZc8qN0523O2956Glux7RhgkQe4ZM7yansHtmJJiw74HLlyOMBSqwa/
Xu+X8rfKch4zOIH17aTfy8iGBH+WiqVXAVcNUg5372HOIyFR3rGuYw+007hCbKF9xeEzBWGirO+n
HM8Hz/opD0jq5rw5EsE9cboYVB1jjjLppiCJ1fAVWjLKprnFe+2o2PWoWPitfz/E9SMuJwGfYBjq
xyr70KpFzUpLc3At8/cFTeiN5Mj5WmQ9deSlVax4rGvH+krjTr8aCbDTFRRSvmdy5HmX7RlHX3Zn
NJdaJX+v3H0loD4r3+jDJWaNdgJPPiQchrHHlfosW+a1/QPTEy4wwuC/ZuSB7Es5quEjT00ibXZG
lEXa28oTiJ9CMUucY9Fu1Q8nyQse/aD3OOPnTk2Om7k1Jzh22SbExfRHJxgF/JLLMNv4fKmJ1ZlP
0QBNSF0rEDRX0PdoXi6pSDA2y1wrcmQ7wuIT28LRjB27PNNp5sVQ51Vx8L1STJ8YKEdeI6hKmxoq
mflGxNFHHo60Lf8HWwBwkLKR5Ezd8hS8oA7dOEgv2BndzY5CBxttzbyPAecP505+7VzmyjXASE73
DEHiwdiwGjKfA2PGw+qXmmEZ1klwJNDbgP2U/x0ahV2Y5ZMJhMeSy1vY5ZUEyMJ0t97iMTfpVq9/
q3oVinrLoQogWx6wbFZtaxLY5wIEph/tWE0e62KGJXPl+1PeSMALoLwDU2++woqJTJySHUQ+IUPy
BuPtgQOVk46qIpDIJf7uWIjBbauZEf3I+ZrNvASzdyPeFwypXCDj7YGo+qgmTfzcAaFJD4vbbMp7
vV1V6mCh9GWFlsBOgdPHrtwsdPmLLoydAOjzjUX/eWuZyad6VtELnqojGmLA0NOrMxoN98Wezw/U
JEtv8ILIxf670idykqGyI/AahKCsx43DqHTAlvbN/19CUhQWiwZPpcmNV2Czut/nHRX4/yGCHhkz
sN8+8kQC2hrKMG/tgqo3AF5Qfmps8dHUBhzUZeZJXmtzKkGvLhZ2MYXbK7pCFeTdhswvoxPd4ERh
NelEMaIkKG3V1Vc92Myfb9AoXfC2+iNav8J4T7Lu+2vcNq7jcBIbe+8EQ54k0NfR+Ap7qKLcrJhK
5d3/0dnclCWWBn9ambC2gtHkAvvqyvwnJthG5PymDEqb8MFhUx6ETrLYAXoHmk8/Xmtel0kTb/5y
l/JmeoY1+zDp98CYrN8dhPzm038iAxK1vDF8zZ2SeLebD+MbaAFlVbOQf3oHb8Eoetc5EiaCXiqp
HG5ET3RkeHsxpj7ESSKxNU3W1BJzB96IP32/oIhgqyjwWKRfCjiP2li1oYxYKCOv7yMF9YGFITe6
vef97U9Foe8ybsOfu9Jl6I2BJfNdHvW3/C707qz2MjKN1hEy5nse5QJVpA7+AxCGaNUAAFT1xWuv
iKpIiW8z62Tty+yReEkQpXExfkOF+/Dle3XbZoVAtzpQLugwkMZKgb1LYfFpi9LFR2EKw7gEps3T
6tUZkRTVQLOjqOJRSEsKJToaGh7oXuJLCXtcApzwJgg525cEfKPELsLY2tsggkgZmCNW+eYRhvks
7fXVZHeR1BO7R1wfF0zGWImAxMrPCMvmjFBB0bNbXQxLFODkcpNqCWRbad7XYnLA1rgpKdcF9d17
SRnW/LZTP5Tz7cr2Yrfrxw8V2zMTGc0/aFrBZM2/vn7R75SczJi8rbysu46jCaQtiIvpSeoYPeI+
pqdV+z8HFNJpsGB5gnbED0DVw6elfGCvp8x3BfD/wKnEIg8T/mzX7K2nZKzJrcSEGO5ILBlMRe5l
rwIGrjdeJSrQPhQBBPM+ttDzqO09SBnD3Yv1/niPhvQq7O0kRLpME+FN5QkhW/UOlZIDfBGCby+M
JsOliZVenvnuMcwbXukD51ZGFvMBm0h6qxAHfPbBU99xfYracDp56kOe3aNnEJAX7ltWpGD/tY4v
Zzzch/wLOOFSB/OCE9HeaS6wJBYZhLC9o7DkqfEJYOC/Hegf04D1Ft1JniSdLq4+XRUxegzUi1Tw
oNSKUwhXqIxdf3wnZGv57eOx1fdm3MaMYDcUuLI5Eb4f3v75jAe4xbvsWh72hlbCbWWfl5/L1vgI
zaoA63KTy593dBEdD+OFs5CVZQIrsu3rpnbI9B74443ltnKLdPjBerp1g6u9yNES/ZCtX1igt9YU
BmOkGLAqKvs/qpjrlIqh3TtWOlhv4gUGb3IeRIWpkM9w4WxNPwN+qOZ0MNV8Am6zxwrIAm26zUve
OPhwi9/AoXVJ/s6+xfrkDvqA7/GdGX3WMxY/NBA/xSFPhfcWoJ/c5ro6h/oD8MnbOBQYgpEqkXxA
EaFuD2JN9cPisdTddsQjkYSID86Z6jtuZVkeKK5afV9Jbgk6wmZj2po1WK/BxT1FkF9YFCnA1Vja
QD51yxNbLfQ5lorX7dLTP9tVJqV9X93iKleLnEG87oxOVeJiC/lGNM9IPg4WUiAu1R9Tt84wcW7T
vgu6DksVyTGliylAXjdbXpFbVFMDDsUaqgV6YAZgW3FNjzW2jJEiJ0PJv2Uh2KS5Em2gFEY5W1ql
omyUDavCyu4suThKXamax20hfI3kkBSvA2ZDjfb9ra76BQkgBOuuG8nKgDeqQ9hMai1u2h7xsGSr
XLb/AxsXYYJTo6UG3WkMeuCGXfrXJiIXemsdPbI1j43Jrcj8J+fjp194kVgLCO42ESBgKWUdklST
7e+43lJHjcH2MinMXyRU4XfXhWqP12SlAT6OwFvVFJ1GtqHK45RyhBD+BoN2g1LRaJGToCRs4qRU
6YQKatAor93h5BCjieZgnQ/xwINhoosOU3Auyt6m8+Xkg1QUqBOUTuV+ZLQ7aYSmaA0AblGKBcRv
iouolGK54WAf+epr3wfB3Ec2OAFoQno114XQCX8pGFEax3ubDoRnITV0yDupCPiJksObqnnT5zr5
spVAISf8x/sJiXUASCY0F21znoA12iTW0jCaV7EbqX3rh7Ty+uKCaBMvJT8f6KoOVwaUG6N6cEQ5
RL3HiV4Gz3PTHW91fs0Fszc0QgbOzfnO9T+AdehewHn+dzYc7zxiQmfE3fKfXWKPqRP2IBo8iRSd
YZHX91Pl7HbsdhQXyYdo1NLEdGbBP8w76zbKRVgLZtATvM7XYRZXw0NcLb9bi8TSbJa9Q0tuzVTx
249+S3ft1AaMuK+7t1PRM08Ae+ZycP+QFlTtGdB7OqSgBswi/drIoxSzupWOm/+whLPQyVqUGslA
CsUidvL6PIgbiLHOVfbW2mnKlO4Ua63GZiXbo9t/A0oCnIXfZUBC4opiUlWAwnAkd/EththO+69Y
7oBxNCbeiV+Y9M4Tb3SRPArn3O7Hml/7t4Vk4CIMPlK3zxJux6xy9k4c3pvi/yA9Yrooro1tJ0I8
tOJEotvuiFIRprOBMsBUy0HbLnBEwqT8I6IfflGhqRngEPpEHJsstPDFxZ98lN872kujPpRYu71s
CMrK3pj/jHolexyOwSOwshIj+rNS30Q00sEPzk/Gzbj+FrZE4ShW+gnWmAeDUa9PWUYKvUgec08w
VQmbXWj8gnc5JNvkgv/c9uB1Ar25vtlOOdeVP4BKvTR7+NCq2CFytsauWZraZesl0TidPVTLt6xV
+9/sxwoP78AHQDMMA7QV2YZLiU1aGaPj0DI6yC2/btVP62CN40DDWeiJqz3TpYWngRY0+PbnzUSv
ND0Ay0jiS9YdeiEeXJLiVEZff4m7pof+oYiu/1m9LCksVdcAirm3x/zbjYqUDGrf7Olu72gSyuCM
1VlcDZAl9Dimx9th3PsJXTLiGzuHeN6yezCXjkPI40NcBQ8YEqF0EpfUsGtSXP1J2ZDZyjZ9lNOv
2oVFeE2FtB8/82+PbqkEGwwc2TY5SDgKp/3NiM0x5X62w17aWRgurxiaVJOdD5fxm/TaNRvtfY6n
fZlth4vocMAc9RmZ306XTuwuYlgGX30LN06sIaYoTNMjt30VmgDJYEqn+o8xr+ny8v79EO170rnc
ywbPn5K7bdP2c0I4nG/s7XBQnhfHeTDb2cekM6K4H93GCeMIU0IlzOZhWOYbfXsXQyuYl8rSD6B8
yzKabhDX5gdqD6eQ7RQ5a8LmYq+IdM5NTtZCTOfwVNipruCXyPimjhZCit9pyzBBrOtAXLaSHrgK
RJjPehDx6C+nximv84UhsFT/i/Lu4mVkGXW2hMH3AOS+QjvfOlPTE52m5CGVzPmoTOqPDTnG59E/
XTdqLHSzQBWeQwF4cI2bAEOHRTSnEKc8aGFDZ5bsZt51AlnoyzBRN+2VSuGo0uWwXTNlw3qzqMla
C1m2GoK+Ts+w/UVlNicTopNjL1dBlwLuFfJvmCupE3m3Ld0c71ZSTEOI1wIaKPGF844N0loIBFQE
CiKlY8zhYn/Txnze/wJ0bsLCdi2Y92F+1gzkFjjdqltjzeP1uSJmsZ+XqxbJn85ga37VAJ5wKsBP
YwDMeZYoyhE4hj4PaFcMYaQW16TEpYLFUzOpCLyM3dXFcPWXGnU7lmwy5StcNzsr10+6ycM+aTvz
2tqbtTPdHr2VzsmFrGdUYsG7SY/JF3jdcQDceordoukG4UW7EcKnwJqN6HFiFYA9KZZycEzgATKe
EiRd8JuuJ+87NOenSrC5D0EfBBaWqRA9umgZKa+QolGZPlo50MAQN+RZDhLzuX4f7dE55M8/eoDB
63QXQvv6xSxPinGkhWtkEnyIDsX07ZddPw4K15dL/QEg1aZVr4B7vNpF5s58N+HL7YW4URSJgL0Y
BHBWwsePtBGSPxywUPmhRKKwAcGa7+6a2w/iYLtPbmzm0ctgfnK8t7FosgygstljBdm/1L/0PVfL
wMAasYzz7JmrAxABP6ao7c79NjOjNH0FVW27faw0IXpBrjf7nGEd81kP8Ukthglx+v9VNuw/usGD
FvQorK6Iq4Kuxz7aVIThIL+oUvVKjh9ekRp4vW6zbGZ3a2VwHmj8f3m0uQTBh7fUbRBqyizhoQB1
+MEn/yeGg1ExVHqv93d4nVsPOyfgXPphdrZ5U7gby0GSTzfZDfbZ5wgiJH3b9U2SWDR6jSVucHPk
lo5p3voWBXVYQ3Skt9P8+oRuGeKUcXhyf2BU+OS41V5A20bcPbLvoYxT+xPi02upFTBzh8oKiEEU
Beh0atU5SHeKn+IX8vluSx9n+G9Cve6y8Vhukhx+X2ETvz+zuNLDVvnui6GKwlavGzLYBPjqU4By
DVuypmIE1C+GEJ4MBzvZwRNUtBYjzKvCC/dpFs+w95minTR9dtqUlRmWU9/RS9Dw6NARrl6Qqslg
IWit+ZSjS5PZ1mxzIQ2CEHXYAHgzPvrjugZsltettBc+QQ6dnChIiw9Tm6/4ngtmoj2ZroMKxrCA
3X1wltsWzxWrzfyi4Ic2WYuv0/SptNUCVT5PNZm47GE254qE0HVTX2VVQoU1UyUjg/a4GnqbFwZ/
WaGmu6GFNUooQVfBI4JoQYoqOxlVBgRZC9kYnvaRLrn0ONh7+K0ri1FaGR9VUBiF7KqD5Krb0tsI
NAEEWPvLBlhw+M7ehpzXAhnyK5XWiRk7NLloeqZQ3gdWsRpzPktlHmDhp8cyF66qiC0Is9Cf3QSN
BjVw2wxxZqlD5SIqRhraI1odUTkAXbq+JU/6yrimCjL9D9g9/EKzGE9Ul6WB3jla1luJisOGEV3w
63wHrzT9rMhDPDN/p8XITMnaqcpRL0eIhEdKTAlf4SHfcUyAZYngrwjj+lojnJM5pLyxyvNVkDZD
GjipRaZMM+DKgYjZrmsJUVkM8VoLNVANrjuhqS6FP4JaV6Qc4m52qktENsc1hJqWLvFu6jBjXSTc
PNE4Q8XVpknnFujWOwFx2GGcff/8eomC4Bhfbjerzu/0qUp/YWQBUhbNj85CeOtg+Ze/QKTXltmO
4VwL1pumDwqQFDoT+kVpyQn+tAMD9U9HlCbjLnPBuswZCP7ze6iyt3kWzd8A4i98Da5Xe6wJ0BRN
HV5V5XxjgrXZ/C/y+3kdo6q5YhT9qfofnZ8j1BwJNKs9CSnkGjkcD44Q8RUWarSUbmxKqeOQVreX
8mnWytmJGw/yeJme5DE1/3ZpJ9MJG0hBD0qu2FcruufvGi+4jZllQF7wfBCLfWgBt31xhq29mKNt
5lXDwZ/UGNcjZcZeVwTdHGUQ4kaq+dK9526haWiV/prOUZoXD2xlCKTEvZT2rS+EoAVIfDGHu2O8
4eLn1ZI8KkY98ovY36A8aWe7/U6stzn4qwc8AJS/w+tLV4cQEuABXa1/lzoiMdznYOVqZCYoZUAg
7GOKxiz1IgY71lZfEJiHTcZivuKqYb+Q/6osrluyjPLEIPKFUch61WSBkVDZ9zmB8w2wxX6otJbh
Uk1b1c5b/6ICUcvgFGbjrdW8CouWYRP7x3Dzf68GYNC4vyWXAwQFme9dwiStn4po8zXwHlZ68pkz
yN7za1VeT3qO2xqlSM1svU/yk5RAbBbNjuZRXOPwkEZIkRYVfYT8NK6cs1jYETS92jcjO41jc7xN
yrBJ7JFc0p3484IjFoZTmyOb3QV+yi+uVxpjVAWgSuOnOTcNfeQzm7S/uBFGtpRxwIK/q5JMdwBM
4Mi8fZnHZfHH9ZBJxokyHDBXI9Q45ds484YqtxVnRnh0OIfI7G2Bhz2L59YKoNZ0JNAFUVnVKK7h
ZAUlCH3ARMk2on3VvoF0uKNDAd02JMqDeAfs4udJFjvKr2mEoGXaxOh0N/al9a1cVQKCCVcrcMni
gh81VvEq8OURtbfdwhekQPXg+0Unu1woXoEl2uVMyo2fx/5E7kkf8cm//aMt9495SCqUJ0GnH5yY
Uyawo+mlOhDVir9LeJDaJqTQUW8Ze8oaOwPAJ6VrsRRpBeFgHanLvAJFgUSZk6pmNLx238V+RwLv
2hW0t/LSmMyJ9bsaf8aKx2+SBj5+qZ3Ts3tMB5chQB0q1pcf+JBae0LiiSIYqxCC5dCDR6IlZ9fr
0GEQFVMZLFPF4ynjmEmHv2jQPMrp7ZlG5EvvO/ny0++KlaHfSzLDDReQv9Dx4o5wbGjfgXg00ebt
aHY6ZGkN92YX1RyH7+JSJguKUZVyH89Y37bYxIxmUSXtzMg79AAg+LfZoqb3o5J7Q07WpVwEoSlu
g+9wXlF1e7OX0+0Z11KpMpduGdaommEBKtfp7cfLAdbhQ8pywmNRpI4zxCuRe1r249Z/FBFXAb7c
wkGr1iIPsILBzRmCCU6O5dFoeyWMdwDlcELR97L8AglfxQYyPoq0zhypnppoLt8brLBZiWOmW7SZ
T8hzpMMpr9qTnRqHeAhs4j78hw0GYmm7P7BcHdujJ/68SnBQs5TeaerAp+EljA3hIBAY4SWvkALD
ssKb8sLiHZGIniCOBnY/aDkU4QgHsjezrmgD+aH3fMddAaXsnSU8IlocM4fxJa8ogkuD9QLpUXc0
aCCzh1RRHbGCpJFLBTCG8Z5zL7QpRsRStkmE3VbK+X/c36OB4cSqvAcGkXmHwFsnyHrRYSCGoHi6
Qg1x97tjp/dm/LtYBEw39R969l2hE5afZE6ILpl0qbdCucc3+fdlwGG8qojaGPFz1+Qu+eXFbwO1
GkR2cbl1wpdmoXsOHMuwXt/Wr0vOtpcqkLWqURn4J28hdpoc+//yE6E8TdkKj51BO9gx/69CX5x4
g6h7x5CblQc7BZ3yV1P73bkM0eN5gxXoyU7K7qpHZHHxFnwzXtWsNp12l0zPUQcC2frL80y3NdoG
otlhSUg09I5tbvieWEpbbnTF4+RFhTFfVJcujfiis9ZLIprru+JgqDp/3BBG92x47vN78BhdCh/p
w1Ii8BIDkJuDihR1Qi4ueDPbIp/ggmPXjS4svHp1O4JynrYuCYfkaeA2lSRs3gT0Tk68fyvwcq4s
PKigSBTjJpvoKZ3HB2Db5sODfXftgv2xWwqzo2j2+Y5l5ScOga+9RQdB4IQqXHSzbGNGQWarQg4p
wZtAVLC1h/QidOj3V0VqhBPZrN3iExSHCm5hFudt5LPlNPNVfg9h2CIf7pOzbXzyME1uG/sztt4N
B3U2XG88Kk75JPWem1VBvpiXarQ3AbzVZInGnsM0TLWTeA+XCzP9OZFcx23sdCSaLQTkJUTiFRG0
MLLZnS2ZUkMOxMiX93lVlgWgh9b6U879SIFdtGtasUk9dcmbB7PX+rYfQPSYOGtyT+cndjkp1IhU
pK91xJgPLc1eFbt92wDxjIyrT3yb0t7ezm8TRbcANHEtjPn8zZkkhZ3Nglky6f9QBDaa33l5CVVk
VOZXuFYmMa+ER7d7E80n60d7jBwYSYsROzvS2CxZFNLsI9kVuHSHqjZi+WiIwQjAU+TMX3B8N40l
kEcWoEsdZMThC/efwUlQIE6xSa4W/yaLxojR7lmLBeHFLgTP8x/YH+tzetL5Uyn6MR2wmhmidhfx
fG+5VGdfDd1eVd5Qg1UCi8B/nctfo/0BLhM8QQQXOEyw39heg3rAT6UXskcJiTAqJ2B5e0ZXRD5a
X324Ejb+N5UvXfp7pdxsiUKQ8ff3wEPT9aaNbz2cunJ+1EQ42qeTjEP3J158wWN3VhcER32LFaxs
1kKwQLkqi+9AIOjYARzmTFKJNAXbHl57MmswoWzKHwlS88j9LHHMKwdnAkDPFOZ+MaCGQMYRDcUw
jzANLA9JqanxqmFF1xe57GbAXyb500Hlq86p+/bPcrAcftfoCGYejFHt88tnxRXlHnxLse+A1+NX
3iduzMFRB4tfYQvBYxwD/AXaqp4Sl0VMp/e/40eQprdhJZA+QK4KdT1vF8ZEyMTzAYR0ff9AQwCL
fHEBcjgxyU11iAeSP1sxohxhxbZa+/QEthqU4fCQApfcpeDEOl5tVviqfu9mOoUQf0gKDZdWsoi4
TxegY8mqGa2D8gnwEiRiRx8WXui0oZgIunVVf7MG9dkUXS/C2KWKwZWrv2Sg7xHHk2vkwL2AZeFW
AOzM0iDQmJDSHuTunfvcY7BAawY1Fnk8ocI85hQIhvrQqYfBAwLd0M3U27E5H25uQo4gLJJLNSAr
86gI0HtQuyFe/2t4Z250baVG9uljOoxN32yOClPdK7kkUeOrPxa18mNNOybPKK8/1X3TIfXJsDV8
xLS2iXUdJaZCzY70npkGKWWlzz/Wz0E802gZmFpTwlVJ0cpNg5lUO3rkkiaHHxiHM1r+nt4AaauK
5GXYgxSlWNlCKYQbAthN89chVlE824YqD+/0n2z2aCUZeDUuAnfvIhTbKML9l59/ijOeSvH8d+FZ
rHBmz3HeF7VamQILxM8h5+r8isB0DyuZECt8su5APw5GiruGhSmzznM1u3RRve1yiLv6PyjEuO0A
tT0jK4WnrLR5grMneSp/wuEnmVJFKuJQ1qe1CXqGikjNOxF+P5F0X0hfxYapKngNb071Deymjqqb
TKjUSH30O1tfyhPsOBFVUuwZgoBIQ+7iytc0Bjzn7qOkkjBjxn9aWTzNIrQit5+xXXCmP7dchgAZ
Ww9dGxI6dfKV86PBBuK+e7FsMrW0GBJ3KqxKHAxlQqTeAmMOE84jFlZhM3FMZtahyhLUDkqYp7K5
FgqUGG7mxk+AVPBwTdb/ac+BHllhDwxv1yRZ2nrUJ2XwKBULQIwyKm4/rG//uIxaAE7c9OWjd/ST
LD+RMlo6yo5mBPLNjNmbzQ4FKSvY0GU9iHhdj/hYVNROp75r1QtacbZ1ilkzzEJaj5/LfHOJEvKA
Z343x1SNoyrvrgyAQortilphOuMZDoxMFXzhZAgmaI/Owam3AqW+WVD3zTKPiy8OmH1iUt8G/mpS
K43w7tYYUbpccTtcAH0NXp5dX4GytpRsTDz9NlcbJ0YzSKslV1b8YA3k/b/2I0d1wZN4WP6/C9lQ
uNmUtZ61v4wMdvW8rCionDe5u0FSQ/8MbIgF6iZ4hUzMn6KhzITBi7OPXr3CB5EmIaMxtzHoJKhf
QbyyBdtdMwPOhDY/Ytf2mp8kTjihd1+XHXjquVkCf5g2HwNduDlCb0h9M1ARaspGJ8Ba9IOYfTHb
vysluhAqcrZmYAyI2qVgManLhFR/rFaTpg8QdYk3l7WhDeAoo3Y5ZfgAsq7AnjOvyOWKh+M8rRDZ
1OYyfWxQyj5hyYTdvXwVCMrsBq6RbeWdHBIPh0nzmBODO0/nh4v5tK2rTL/trLyi/CUYO9JQYT73
CgFpz5MFEs7JZWg3CwzIZKjmU5zmHJEW5SxIWna5Lx6nLNnyyAD8jkW6ycDM1d15QFqsSZN6jjIG
0UanzllbX1lkDKMMUQrhicx51LXlYchVnz75Xx//OK1/mHcnOUOuJd94NxrWNc+Onjul4sABmjy2
AdDtjbuzexgt6XwKeMVmJkRLodAVWI+3cfKh/2s2WRpnPqVJ7DmyqVLQs2K5oPveCylHPywkWoRX
+3uxWtKMFhtSS/ufnqcpGXNN8QpbAaW3PPlA+MulDNLhzLtEeSW3dawUk/NMWC/E1ajMQWItEIdc
UbfJxyPO7H4W5PKRJizMoLz1O3riEwDrVydf78/yuZW6kl/c/qPUqjUAiGCLDWlYUTk3S3X9N4YH
Tg7MLRJTbMan4nbS0Ysni4ZW9xocvm2qhHVuOTnsbRgaC6I0RONvn47skZWK3yVTTv0YYXUzjjHx
6urc9owpFCZXRsUPWkokPW5t7WmWtCly6NEC6O1CIPM6O1Bmynj1Tj4ddAyCPgQL1GZxfxMbiy3t
ofEhLptGfj0uihyh329qmBOTsYfquDn7yQpLKyRlzyIMsemugCrRjzhMctRpxWVAmWy6Gy599G9G
HfcN8VsCxsWuDG4VYXSZD4GyC8tTDYEb7O1WiYv+tPv5AWwEs2TDt8OnwrLFUQb82Y3vBFtJmkgQ
xcybaM/3FJDWMVWe0Ka0GaFKxSnWhy4G9MLpHxZZekPwCTfAmBQrxETNCUipM6k0M8ZCqyS/PmgM
Ee5fZA2u/N+DjB0J3G0bGCPCE0ITCrWyQPtMpddpErz48KJY/Dzm4jEwteJYU3qjdh3SAu+Ac2jk
ozTXN3jldAwOUVsZ+jrSQBUOJHUeFfXA30kcSNr0IfpTBBjquPuDNXXYFaeBb4Xph5q1sJu/I34r
av/aYQpdy8Z2Udu4zMVV2DPxJNqr0yKhCGeFVThsLYTvfMlvHuqP2XAH2OVZZpoUBnoA5++YhaT3
DUHgIkgFkOwtXg6oHvPIFlPFsWT2WpZrZkspY3C5oaIzkPus7k1oSY2Hv0I67PKwRTOHXftP4Mu+
W0wJzUuyMh74cmd5YR6aP6zq/JRExonNiv63IDOL95HY2TqIvv+Oy/Tel3/marGKIPMHU5B8zF9P
WPB7FW2Gyxaa1cQ042NdtVoay/niEuT8YogPB/4uEwO2oywfRY1cT2A6j4WjTYzLixXmDL+dU1kz
FK5LmZv0mY5fEx+uxQSuOCSW4wBIoYhDxlbvUr4ude6Vdjg+hlS4Lq86vIv32rCHAvZ1OfgeBZfA
WAo/GsiB0+I3ncHx4NI3jK24r7bltCbQ1QfD7FBLJ3gUhlUnSd9ObCar4uu1/Mo5/bIaVITxLvIE
3slvwxpfHW++aVM2Nynd547GLoIwKP0UJNt/7Sa6q2rnUJDEXdBFKDiaRgXe5Yx1fi7Jj08mzCq1
7KYe2b3SQmjLsmeg1IXC1eqBz4LPot8BxYHEIKGD7KNQHoacyVvcjbzdlxKeyH6A057PwiXAyxLO
S8F0PrUEnZvQgwUfrnuyGSwNeVPM99VMlAU/i5G19uJwGXt3faivOwEad3kkJ0dXyG3toGqs9qz5
mN4PzBP09pamjhff3UJBO1fXJsrx6xWDZ/XIkq6loQx+gJ9P02k535FdX57R7DWlVu7DgK4+a4Ko
ANsokITTViixPjkxImJ31Ojz1cw5i/U2mJitgHIkiPU7aCJeq/tYmKiDmdTI6Ajsqi0+PbaugRjM
d9qz4wihAaCAALckLqFMHu9nbnTlVAukcBXaAe3HR3xabufDKjAeyaEKut1ZNLuEiJ/cJdoN7NwU
rXGvj8JWK2abCbko7sMj9TziG7jD9di89xEH5dLFQVmYIl8qoUZTsEUqbuuszvpNy04YFLQK9FY+
X3TOWer4raNJcGTFuCPmnfflrY9HAxkly1UAiTZ50zHOnAymupQniZPmPHVvn39bgH+Ej+Nt4Vxu
WgnXuUZ70ewJMhRXo4n1RtPWNwHVmGfE1c6lBph+CWZ/dqfRlKGUtrloWOyM76R0KVb/yr+dm4CI
eVyu8I+pT3HlclxAvZ3gHo4WgLL47ABSmpWtGOWLQ2912QOjktPuQPM/8o9b+mjMy7w4gyOLioz0
oHwH9cnIraOLFZtZ48Oo8o/g8gZGL2bI5eB5FvbjNvPsX/w28KgSo8AzMF4D4qgQVcsa4YRczhev
0bRBFRgG5yDycBYw7zFvcUWVyNn6IgdISZ1FnmWTcCA0nMoCFSNM1WBgghlAIgiqdyqjpXx6AJIe
arjv8AWe39OOAAQ3E/R5vPTeZdyUEPVYfT4RieDp7DFyPWY1zoz01Xl3hMCus6aWNQ+GXD3+41zu
a/F0yo6hPGOB9FdAtPN2SZyljttFjjYfs6UZrVk58HAMqQw24s0FcBhEpoWbANdyrKkTHsCkT0P4
sxGCJgAl4GhJt/3EHw40sOg1iwpVxQanLweWOak5uLssVtN6c2EAL/MFedcDFDR9T3Dz4Pe68ItN
8BxdE9oKXgiFSqRTgfFo621X2ihYdbKCAxgG9VKIjcG0SSEZ9asFegZyjzHWhJFstfMzZOHw29/z
G96Pb37zb1uVtowWLHGSJBnw3I8TONQhyZPV055AQfBt94wMC1BAr4p93kSX95gk2AO9/2o5uL7o
A+zfARLsgvq/dxSzSS9j3ktqZBHllcaWn8sYnEaUzdOqJNE/P0Ci/tS4Vk48/BB3W4N7mMduJb2p
UM30ySIs5DHF8GczNVWQ1KAuuBJzZtu/Co6C/FX1PvlRPoeDwLfz1pPbqjLOUanAvN24bbshS6+m
k4oqDucw0pKxAbr5fxIUObNHyMr8Exnx83v7ZjiL36C26sGU9Io/ypO47SmURehABl+lephHkLo2
f4dbhiRG48QUyRzAy5Z6A/5TlMim6A5AGFAgqpsQkQzBAW9rpa+DqKqfVUt6E0RNktYziY2tLxVb
UqwTNAoIB6gZpV1UsOHuME5y/CCs+IRAtpKvo+ptR24gVfZD/p4OApI/44h0L+sYXcHxpx/KhLO2
sKt6x+Q4wuKumxClac64txvacoevZsbe+i5LiJUS+LqN7iyLLN47IyBWDC/9eJ1w2M4JEGYqL9PW
zUVgKN9rE4vkPVYrIVnaaOL1GOv4B4hMqe5+Fj3aUlGrf/31ZhtP2PHwDNkAHBqt3o1Cw68PvJPk
wxdDkNI0/J72NsO9ZzUJoH8Qs3iMbnWl2v0tzElRk9TAVj0gNQRCxZsgHZrNZHAQT7hu5a26CTm/
5LWm6WJJtNMhoaNFgDC3BjYWHxAHA/cVyyF4Vm7fM4Yi1npC+TV+HSJWMWTuG0XGB2L48d5WRfex
HzIP4PkUQmNs+ZvMY0c/VvxEkXEHQhBNNAEcPShVFjEJ5LOjJo/gUFvvoSLD0CylaXieWkSlx2io
xvwfJKCHAup1gMxejKyc9tBxVe4McJ73iM8G/Q+N0m2ZX32HxNRXXNXFr4dITCEFbbXknPIyZPhH
zJ34uAACmSn3SEZIM2eu8iuew1ff4nE1HhHMk4lNHLvcaLH9PuBmxdbgXXBknnNYHKi3JljluM9V
qNTGgPqbXnEyYfsdYIt5l15o5ZbsjBJ/HXsdfxE9EEdxIJSLKhztmwfCN0Tkfxpnd8iDe5kGm8uL
hxCjlzKdhng++lte3v5eWgp25QfBSEYX9i0zuHxb0u2X1eT+B5PfhY3Vqi2G9AzqTXyYQwXzQjKk
cbge/1EzOqZFufMRNN6sNLa1Wa5pIkfT4pzTYDe2iyGlUHMQIEin60UbonIPG/aJ7nr27BqeJasm
p1hghmBgB9yfSGKANOzouzSRstTWSodHAYsU0PDue/BC7HCPF28iThK5msg0p/q2/9ABXdLmX9AU
uiQPBI4dZ6JKsZpBFsJvjygoS5A2FT3T2hibLjTEDDLm4ucL5irKfgQHK/n4LitQMO4qUUJ2fjs4
rxV2o2AdLRuumTwbOEgGKI+MyRjJFUmo0KXFlpXJ/CLzIo03/3nYa03LwjPAshwRtbVXRGBFLs1F
TDWvv3h3f/oBt0xkciSnkl2YB3V1fT/3YRGb14lhfILuYyhvovrTgCFuW4AHr+LfeoJKVp3TVrKc
0ITO/KhxO2knO8R2UEYvFZXDek59+GxahlDEs5/wr4xpBKTdGueMDsLtTTsKBN6PbLYGcNfN0k54
NymYW6FzPM0zuZjmLTuFOzWQWUpl6r1uMwxK4FIJwd3l23k6IwmD0UmaoOvduOsGvt5MYeSK55JI
b0ARJLXanWbY2VSAPXviP4/3YJ5zM3m+o419eBjXnihvkcgj5/b+ILbRJAe0JuE9Foh1z5co3Coi
EWEu61prPWWVlrds0kLDVnLAhj13mKvoV0dgp1clDLbvxbkGjSXc+rFNYG7ZeGY+A83BKfw6+uia
UKRkx6lapl/TFDSj8KParu3C6ZitJIifrk2VL+tyNDXU0KNKuhpqDXjy+cV4TPrxt9C0FRCHXJup
hFPCG1yh23NH0LFVricWaFhGGVB9zPhxMQrtRBo7ALFL0AyYJJiKhXZE9LO5bZ+x045lw7wJfyD5
Ykg7A4VUJgnbMSNf7+o1RbszWZ+lz0k73M/WrDFhVkOPBVfBxZRDIzPISOss1f7EExqT+XHgJbLc
OmuiFaCBkBTGGHpeIoXdYK7+OQmA7DI8NDMuXQ7df5jApvFnQpZVr136IFQYB0jAkVdJqce4XcNG
70ujzB+sv1Mso8XkQWcPl9+0cilN++9Xkxyhhoj78woOnUCbNmmWb8UpeZIh7J9Xst5NUduTUWR2
PgApBWMgI+VODY7akIxU6a5MW/4Kgmkw52QRG0H5T6HgFHqqE7gikEZbhg0EwdKLKNmJV5MEWNeb
p8C/T65MLM0tOqVws1Hb6a+k05EGF3Jb5aUGLMnEf2i2AkL/ydkATguhuqF4SGltnfQdyx9lSARq
rn4QGuKDltMsivKwRYXimds19uC6vd3Ra4ma4bmbZKdw4VFqnLarYPt5boUv15I5I22AvFRHs0uF
4c7K/rZ0s1XTDaoFGmWnV8WfqX3n8fas1ALHD/lCaHvS5MRuQ64nG4RPlZlHomoNxVNfy7BcEKRX
i2ZMgbut7E4RxRHPk2bV6RP+WGGb3LwbzVzZYoEd4sHMxVmv0KHHOMw3odVYVod6ujal1KI7hB4N
SvrwOBqZqAOn6ttDyvdC22bJwiSqLaVOmWkAPj9KraNCnMr7TD+KSoVz7KeOu/leZbHGpYB58BbT
g3S9BBk4QCPnXWfrqTCdN4MLfz0qEIDN8IPcX9yPa4gtNJ0GLSrzCF05y0mEBtyrwN9WSoXUvXto
fPS/75zHZqEjM0YRuPFufSy9rKm/oSgKSV3ML67TfW9An8A5bokAf6AsTd/IpSYEoPhKWUdZRLMB
PxW41aOGFhTEqIInkVSzmZKPV/Tuz1WKFtt/S9I0JDwUMtQ9GxA0Kk7m937PCJ06Ce8QjiUm3oA4
oOuVfWNzaYvFJkjhERYW2+i6emd9XURPL3G49tdZknsgqAzVZ5GavKJYYeCFS+jVWwt5Dj6j7XxW
+jNrl9CCyAjzfQzVTGou3GizSxHzfCasXOX+vdHG3vHskDHmK2+0edlQn3rp7y0B8XkBeQwruwbd
6LYhW+n8H0r5omdtgQ2gUJK+Lgh6lVyfyf9PlgjrpyiYy9mYXNcO5Xjs1qGeGzaU9hFEYmCYC7ly
XMqXYh2LoKSEswJIEQBKZ0fAB/CznJeNewqssEPepU+73G1KplGubUg1b9YRvZNkKkfUP0R8Vud0
31moVhjhQga6S39cfw9k6oY2qZCFJVe86FQNQHzQeR2y/T2WSpQcRJqX4HbXxHI2LuotVXVNS6wF
kUeWZVcElZ+ibDsNmOWM79POxXd2gHhi9eN94VdCLue3gAzMvDR3nVkQ1BPMXs0xmy6LY/5xC1rC
d1pwIhuLBqtkcyIAExm7we8ZMHA/jCCYkSYGkDtYSa0fbwEJ5Q4ydkLQCbTXC4RnTR0oCphpSW5T
/yyI1wbwA6HdzLj+Lt11+y1E7RF62Q7mysDtzp2UR4suqHKfAaPwijkT/JALXJ7VBbjBZdDYi2mR
6EWnsJPbD/jqdVKlPWESOc/qIrqeYQIzwjgB1jegjLzGvwgZs9JuvuW4i5YRxTP+nb7IV9eDaFVJ
Z/zpsXwzd6rhQzEAMhGrOIHeQ7ibZevuaFiVsui60A2T9UQaUn7GB3KVDma1VLXuHPHZND1EdyDc
JBf1H04TgkUF5DKqTQ3vPx7W1xkbrV/PTGUZKPyoBg6hZ7YUea89T6AvUHkAowKiRhvWN/BeGABf
BoEwwaRAaVQ0NhpKfxm848OilcyguJiH15UaFyCCVGLkDbsG7XoUseXV8s39ix2z7Uu0WYdNeAIB
rZKJumDcxaH5A4k+Fx2SS/nwO/dYM+Qk0ZyVo2qZ1e8skNjktejhJgwRDnbcWhMRyoWd7bU03B7k
sQ0FRQb/XC2ucMJlOrf79kd/AjH93HTB9PSOBjDH3WwfVd3WNO+sok3U8KqmczUYC66PqqC6j9Pz
//0azClXNX7pDXLoqcI12EzCIyg4Lvrk2O/kpjwFh50wb5gUii80j7B720ZgEFUaGnM8ICdLaUqk
1qY26Usxu5Xr21oDgdR6WYtC90VAnht+FxUhTvUdY3DexB4BdC2QsLpt1E1SOUUlwD4u6aPIgZFR
5n9RHfOacSpTCD+Vg9Xo9jn2rE71HchAKi/qIrA7HDdRq5V4pM5/2Rf4goRgEjXA02xoR1NxVoFT
l9UvuobPF7RD0BhftX138bKnobHm8BIJK0zBMoRkSEA5o6ocsmbKfxcqg6+nVcsh8L/xlG2zxl77
TokJ+6lBxEYVQbXPpHAdgsgFpcUlTFzUqv3IG8XpX/jDoDUsxKmHe6GH2uBoGO0JN3oUthxGIIAF
R5S6FE3+Nkqm2A1Nfyu46HCSol9faVF1fELQ4lXJMrnOIZ2AMC+EcqbW42SGwmzQicn4qzKvia3V
G6CJz5qawmBs8OpnWS8RbbqHVt/+t5sgnXpA0AaD3D90+ao4ZRYJPnuoIfjQ+5ZGiNG5d5F9EUn2
RaJ/VKZUzNMwJwnWqt0Wajz+eI8GubWSeUV+X1NmzjCvmjWx65O0bbI/cOxjV20iulvT8e/sJxjT
qw77rm3PK3ssAcp1KOSEBOPnPKi2s+NVwysSNww7ZzhXEsRqYgtG4yADtpy2mYC4rkkBYLLotVB7
2rv0Kln4eW3ApyAdWf83CKmCEDoe5fU4DMZCRTeRsryTp2dXKpIleWwfjBqO+nGi9uQ6KSHAOxY8
5NNoQgUp/kUiEvHCkfL//nC6ApDJMgrOtoYzvWoRjbMBz5yuh1SpZQEpUzIzqjZL29RncJnCv/Xo
Ug9ZUv4ggV6mZPEKa62aQ9I2CTejdMAyDw4zW6/r4TaB5genM/iXaIcIXVpnbMw/RqlySuGOywcb
7UhocEwu0FVVAtiUj++k/nFTOcxRUtyv3lhIx4/bSdt+Xha4FKvP00s16OmShS+N12lgjo3Bnz0K
hbOSJSQdu3fxRt68sz2+NoUWvxKhNHSlQejyKZ4KqZLSjyPuGiqPbDLhDXSX8I7tr+0wfeOsVPzv
fOSYNEfpCbyYlL0s54+h/kG1LyeAn9p+lYmU8B4aGYExSaTBa8jZXjF5BbBkLqoW6hJZjPPguZSH
SUiN+LFmX/rTgnRnt3Nj8mfO0q4fmITaJ35S20dsXU9hDOR8cwn0zz3FYh0aX4sDdVkmoBp7UL9A
HgNBO2KPEoyPWIRQfhs6g9FE0S9gtEun9I5tSYhqFiRIROOkZUxtCfVZ6Ohyl7E6cntR+zM4k17b
d1/dhDIiwEFSLTR2xhuUISK4pmF2TfdEGMZ5Q5mD3rKdkNwEty+LzsA4m8IuA+SQuay4ZHH1ri5O
4mVHBsgAemauDf6qfQxbgkng4zXIpF31wm8nluUpA/Pm+V1mWvdqyMUCXeWyp+WQTwLxbCod+u6M
PEXeMukgGv1z9hx6t8Q4R2JpkDIYPRei1OW4xQS71fvOKGzeP/rPOkIsPW8+2sJZ5ynZ3kXQTv3v
ULw+TbHlRM6XEBSu8Ht3AiH7Aa5oEVaRAp8xmoS1oD4VM5xmnN3sCasFZ2y8FU9mP/j0Qqrq37Zb
qytFXP0OkhTDrvV4Qg3t/VBOPV3iYs451Q2sOC2MaErCz4vV7aV8An1FKr6upSPJD1WuM1VKnf9s
G0bTs8Qmrk5Scv7A0ksQCL8sVgY4oBPc1Pm4sXgY8LH3w2Ra7cIa01ldinbq1krKkdKdYokypCVu
WAvRoOblkVW9tjFmsBcER1zwOsH6mQ2uP2vq8OHNFUvbN4Yc1Wf9O2xglF4+Lo9Qttjdb5J18OSM
zAc/zYOOeBKJ/8hz+jdMeY9lprxRWBUH9UGCy2wAFrGfAjPms6Ndxpk9oodaOUQf6329KG9JG6Hp
CR71eAqUDcVqmuj5AqVi/ImNrueHGX2N5YYtlQKtn7zOQ5xikAgQW3ysYl8PY7FFbUA3r5GhWHeJ
cNZu3PwkQkHog+3R/b3oL4I3i6G/0dbkzqiQddI5v17yPYcrh01lcyLaNOPxroIV1v9zXIghS9/u
WPKs5NmDtOmDdGD7QS8JadnwGzwZXoi2WLO0Z2sCzpNRq/Jw4xidkt8qU7weg7CvFELKgb4BNFCn
idLyqCKS5OH/BHVulVKbPi+QSK5ERhrODXA97kqYOFeu++WqImzYk+hNiPCkJNJVFADs4bfhu7Da
NLVP0HdcdXz8HHL6TidC/PTmmfYX4QxC5HYZKIr23OpwxU2IRezVO5l2AVELIFdTcNwyqMbLbKoM
GgG6fZNQG4/OLhu+u7FW+w/SNNJXl5PL9/MrHHgoVQX7yCFeb2D+I5pwev6EdIHQ2U2GSIPs8XT/
6qXV7fwta2LvGh8zeSRFy5ygYFEKDEsLnzSUfM+spHFzQu3CpeKA2Mw9cyma/0aIp3tczfqGeuu9
UWgE1GH6jePpP7u57hEilzIjcLG8OzfquXBecUMFC3lSgAHZ0Ljlxh/Q65YON2mUTRVu8q8PfYBo
O9lXb33nucStvCkrJfqSlqbFNQMXXqrKItI7sk27CDeBMrqxLT+k6wM7XXmXaZVECbTtDt+cxNrQ
1B0itDo3rVRM7Krp9mCqxj0RVG6nhQEOKocGOJXEdoMv+bRQYi+TAi9hiDsuVkzIkkNvhoeazOgk
xZgfSTspHuj8G3+kv1KDVTuaaq3QV8JoLkKfVDNilHy8pzMMRLub2q/i7ZbvPUMaO9GKTpMQ3s46
Df/XSCNUc9FKFfsz/rbbEJs4CbYpXBcvtG016M4OJzPeiJU96FzZPulXZpYLUMnyryuNGA9YmYe0
ZDXoQRn6S4AAfT1USSlG7LIWhXLl8dMIlXtj4A/UE/PSLZrKAJgOrn112XE0/67R4ByK8knKD/UY
CVuQSl6ytVoEC/26mlTTCXoRI9LQVYJuYvUkv37XDGbsKhjs/pk1kBrgSY5mDbkgBejUnCX1/Bsc
KAefuvYgTv6L+lE1AINPonl9+9UI+7JHaGKkS9cdXN6L1E2RhMIyihnslf8XYIsE/bWS6w7YKuLy
ZXCU4Gpum4Q38iF01t93m/eNEKWqgZjI66j1zcMMzouovhj5H/tpeTzjZQ+Ka1ReP+bgoGa07eaC
PBje6dmXPu6SZR1VxTKYU3o9Dnfxc+IN2Fg1mTHHyMXTc+pNbzflAPZfQ1oRHpM+BDywjT4LkM3x
1BaI8A4qhwBaPA6+2WEA3NO96JRiZwLcJMMHBpZ3L/yOsuIK8id8ZFtEBsVphyACM8OAPbqsPq8i
kJHbsnSTPhargQTjhrI/e9Hq1K8Miek2LDgKx6/H/ph8p7jdBP8DaNmLPXILBd3/QUYBLkSmm7Ou
r3U7ZIW5JM5kQSjaisOrCTUdAOSrj6B4p+QdmgGLYutSRaNe1oTGZL6UKbMtCu2346m2Z9M97fWT
9Mx5FFdkq9wij/19j5Pov8DG05NgpiU3qgky8QQLzinYp76HkkeMOnRg6eBLuwo/YAufXGPpUfk8
ZU72pvkKk33zCRyZpBe5t/PKwoaO8ItTkLYMwiwU+8F3I2oKQ342f2EUg9/EB6vefztKx6/Cjkpr
VNge5nfcxcTAlk0zfx9T+5k+vOSjX9lfvbdcZgbXqDIcnHJwhZoS2ueTQbT75K9n07AosYlxy46m
eaAt/t+e/yXRuSgoQUJq37+Nvphxif63P0pkdEBsuSvlSU2TPBRceS7ObeiHnBeiPeKkGByovI7D
r4xfEaW8efwKZ/unepEfdjbYujwkD33IzSkENACkxIn8gZljLzQdTU7UMLQ89DfshTWplB/DtrUT
hZQ5qwIwEWA3pT65/nt1LzWXjUjYvURZUd2sBbM7j0UoemXELU/uNBZ/sriOm+nC5V6OrC6N22vU
6zYVOBoZvvKiC4t6n+dbLYidXec3QTavFPIGvJGcgF6LF/Ia9upOTW6guBhSYLmQEbPfhsmjF7TB
zPr5CiFQVLVo/f3hPy5W619q0epjhEksbqwmeNtstVJdmf9GTAdVpwrh39Ks9ySHcDE3eO6QDNDZ
gVgLkjye6/h3jBz9BVH1Y9W2/M9eS8CPqwKv9HPGJuIo1Kz+09kmwFHIQiVK8P/TkE/Vi9AloOKN
1w7lhMJybFtpmPM9IvqWbfcOqgnGHrrfmr0XP+E6KF/s9X2uqlMz9mWlTIKm9orKLCOF3SabaOjt
tcfsQFhj61BsBuxYrbqY38QTQ4Su01y2qQMWwTwupj9auFH/W7PYTT+Fsp02gxSQpofSrF1UHNUJ
J87HMb32kaqi5/2KwF7VrS7YNX+IiC8pdVk5M9/p56M5CyqquxcsYTdE7G2GVlelvNe3bgwtLhCl
UROiQySKbY/rfQqgqkGHkXqXIqzxIlqnFc6A/CHzDafBMQRq2xJk+LbyaTwCWoZwlbT3BfoBvxzN
J13hc/e4coVjn3HfHLruGVPHUXlZhsynA0OAHX1lEFkS6KX5hMj7FT8h/E8JRPxHYNi9m+Zx+D8D
1ylpVFGWWCUM55JEgo1wozLxw/M5GgmEazjdxg/iwYLmdgFgsUA8pDJTQw8JEW3D5BRjXDZGxHbv
6utTr0FwOuEUq4Vt0HqI26ogwWltVJuWs8TlZS20OalGS/LFbxQnnJrpDYWN5IYm+HLORPj/iYiC
nQby+yzuDdcp+ZKjI9+eUAXf83ZP88n8G8GiylMjkod5X461Xol00BsTQg/j2Cs7sr3ZVlhqtggK
RbKPrLVzt46VGSGDeVML5oTTgBNFBRPhWaDq0sZzTmKBlSZ8xSM7jKfh9x5Y1qqnzgk39cehwKLS
ikR4oWYYeseW4qdpXdmxy9US+00MrDvBEIlToB+KMiPV+B+kHAgKBJoatqLv95cto08IiESohNxf
t0/5yI96FFdHug5Uy0KS56MB0pxudvE//8qCmqmPMqJcQ/V8DuoCJNiPoNb0jWya/CGyNi8OPF+P
W5jhZ6DLOTRWRqyMfZA9USonKhWgh9z8hejAi1PW+1pTyyqrzqcAuUBq4EKRKGS8xKrjKskE2bMU
7TdJAqd0kW2wLQ13Ree7llBoBAgGHfQ+vT1BDuvlddjsZYaxPedkRm45/UwDqQjoiXljatS6dWM8
E5OTAhYSD4Tvlva3uXNRczg5bCFck8makJSAuacqHq5EmYmB3lU6eaJqnj47gt4hoiXbFe4s6Z/O
hETEabfGS07wby1ERtS1F9Nv7w6G851+OwZg9/iHISca/f6WIGBrqEVvxu2e/VgJ7oz8zP0Ir+AS
7NMbBJLoxSj31OpvkpRhBwMG2YQali60r6XlD/88bD6XoDIdNHVtmwtHwHAFVsstbtMPAnuHmmHV
D8NkN+z6qaHCNT5glMktbIcTzDX/aKT9kkQphG9Nzlbv6O13D3eQ6kC2n1oQSkacdUbIwtk/ZxAn
YGKpqX7A8umuhGoF7SbZPDRy1xVh/PKpAMuscgXcdRbOk3V80J6jzXz38qx7HiJtvv0pXzD+66Fk
v+y2Upls4MQ6JswUcAsrQpkQoUQNuNW+Y3bcmntEHdzacoVQhHn4yUj4HcVHdf7wKpxDWkhosI9O
r0PgT7L8I/GsVhVpzIsHnJCR/qdzrgQi82rChSihIqUtEco3zAon8NSPcObT6RM6L6NH3ksKcblr
As/Qj12t7cdex7dR7urRnFIjIW2C8KngR6V2nYCrM9cP2nd5gNAktexSckzHW/jINDCIlGftFMdr
MKs1kRpRbv9zzOvs6cZEluYeZ+AjTe6ttTmfbWpwsWGP5OUbeIAq37Xtmad17VYC9KZ1/PWc0Hjq
cnMqSD+qTWD35NLaqA/1eSTm8dvxNPjOK+XNr0DRUi1V8xzIzgiZw791dx8vkIwiBz2ND2sBQOkZ
luGeAa9klw+HkSTuaylezf4S6C8oNjlqgI2o86ZEQtBiJztPThJXFU56W6qfVDT4utGYVRmjMWkX
mlBOmShGRMMiTyPZzWvt3atWTBs1SWYw2I4pnOnqdBgOMtmeROFgl1PqsNWv4FdzUPRUAtvlzqSw
I+PNcRqJQ3zoEPxmxifzuLI3G+TmJN/tgpfQ1t3RfQlXia89HhilUdWl+m1KwJnec47lgvfcQXVC
mCcK7B07NonT3UyqnqPJQXxlIWOtp9kX/dV1mYOZk4hS+Y8OZaMMqufJYj92UD5oaov4HqzSs5H5
gXNDO+6LVKQtq6IBnRnxrs3A+hteSxuulArqWvX33ZoD9jj5uU2zi61rGVhy2SdONQbZdESkloBz
Z6mgoKK/hn2eBL2q1j1IiSPldwtBG7ASsVoM71iEYG0jq0b5nFtGwm2MWSpYSSBH2giimrfzYY5s
pdtzLgEF35rlSYnGvDh4uVtlyF0k0dZK4UDWXFiQD/QR+5MgYqli1D74DMtIh1szOvRFZwLzBQvi
8QwQaB9W7ZEa5Uxs16RrgvYTzivxVAozaRWOtv9XZdCQpCxVQDUmXocU6Vx8M9EZtPwJ8pLnUDkm
HTwWw0teCVjv69SLL1GrJ2VGIkwajDeNWDV5yvEssa7G4+9xVZ+ALfrKd5+9xQPF1XECGDZfGEE2
AZjSO3x0Ya5Sdq49zRP8uxnAiMBB4L1Ap3wCMLJpELPSqyz4aedCc5RJhD0OWBLT4Bjp+FD78P82
cflqPfLFqwWLJGyhkf2vzdj1SKnYjqw9f7E0DqcYIoyajZpfzJVXc8lNQItkd0Bbivh8nGJNB2Df
wjyzAhzWUU6ZbMY43A3tneAOVHbZ7o2aOtekcbfeHIjEZ0ICAPi2MFE4+JgBSh4UqE1A4Uhm2XTt
rfCBN0xeNxiVZycjmOpLnpGpd1fdzQQ+5wgOFPzvLJIbhKWhuovLNuo08HcChSHjlPtfiG/WhOSU
Q8DB8wZNmn+W43YMVsLmP1Tzlc7YphICLCHhXMYzpuIj7Fb2AjPTg1MlX/ht63fNZaGyCSuVXyX8
1Sg+koMJjvfXNrPTfA2GFyKIV3E2uRzvRBPSJpgDZhbaPvlYO2/M12Q5qMl8EPqJPl4sl68//Huf
vArym9f31Bxw4RwtTbN0R+4/XC/JzNAw8Z8d576vzDGsjar8wAxOgKwmZ54wJXzJGzIgWi0UaCzZ
AwvzjwLk3TEqmTzTe9DUQUTriR8Anq3iXKPGiLZv6TcHVnIL3Qhdejvk6lhlCMcBFI8XcIezRv2s
Wm+OwauxCmN9G8u6ZgY/3mWwK40feltwHN5uK8NgA97yR8+OjfQekAIXGzGAy8NH0xCbJQqSmxw3
9tJbG2B+0mss6lGhCgWT77Mveji7Tw+nyJSqhFVF/u6RPhH55brx1ycKpFV81JSKJlOwIFVNGOP6
R8aGbZq9hoUHbp3i6fywyLjSltEBGSgeqi7pPNj2q5UsUNHdrn+d2qfFf/1yxBjTB1Fu4YjZRphP
ECd71bPaBa3GpaMx9BHZD3q1FYYNtVosf+AgyQa/lo7ZvKn/glkE5oWVm9RbPRtCAfR1asXorIfB
bzcFKgldz1UE29g4Qi3ROJJyn00DFJ0deOJB/FdEbc5CvgUXc0EP3Hc8erOLyTplUXTpHWdF3RZl
euKG2Qt560ADn/2L/ViZKKF1GC1pa4oZXPcJACrxw6qu2+FMmW79LhtZsjqQ2oSM4LpFGcALY+1i
uaxb0d6iDQUAYBVB86q/Hkgo3nzYZ+z/zqT2N1Fq15LE82WavNxddbztg4lryaS/axWqvB7NojWz
OBgOljEB3ZjZPfiIFMpJTerPdx21IgZyz3xnZD9DKNmJ+IE2XwWlhOcD/6tNPyc/uyJ2IgiSJG/q
7mugZNf8Go92N0phkZOHueE3aHj8UcZwQO7z3NZ77t7SApxZYi+FzuI+pnQ7t7PIoBHztAcgtOv/
1ilqoWnXhaucbKibS/Fb5OOmYZ/gQAlt1o6YrZ/HD8baJM1FgrB3oKbtc5s5+xkOLNPy9oX1p/3x
KxctXqIsbCLuyvNBJiVjx6jLAZ0dH4FG0rmVLMM1KT0fvTV+impSL8t0KuLmrE/n61dDmtMdSUUR
nQxAp2fK6vbIOGPQ/kLtSAvqLB2LHGj3aBTxQ/lVeuvrMMoBDq+n7zCzeRYnGNAxaR0Nzidm1Nl/
mSd5AfgpdEmvVyYc9YxFmCK2gwJy+or6adGZCM9ec0AbBYYwwUzGFZg6gTahuFr4mrnMfM/RLpfx
x2ox6Xb22mBTNN8obr586QfUN4CtPwelVCuJi+6IYC8kemktjjvikGwNsgEri9KSlkZWJ8GCy60Y
EfX1XB1uXr0Wr5YWixkTeUBcGXRVZGMvoPnJArpikGSSFCZH/qUsaAV3r8RZZ+i6W/ymReVFBm/c
+Y9KM8QMwDsE3cowZyUFYeQnOGSjr7hKOGLruDT0c4ttqJIsfN3c5l9VfPvjMwcFF70j4elUVvWg
YU3buGO3IAU8epIQgGaJ4DpayX2ldrAknp47gS1Acqccj7AS37ZLIpB1fhEp6HGuFqp4RBsokvhf
8LAlXlp+wT/EgclzV/Jk9yiygbaEgaHUjfWCOh0sIG5shJRIRFnP+4zSKGaHpKrlfEP4SEFqzHvK
a8rBnIDboc7QybrE86xfaCuZLR4hw3x64ZCYOCQAMlVpQb+Y6KLiyta+kfjF1iC0aMQSDHfQtI+L
/RxL1I3VTybVp8sd9H0e+dVVo4QG8Mit18/XWiRGvg5trBlqAJvfF9W6NGNfpmP7nS6GhOFXkVrk
guD50p0/kLuLXedlcNSs0mEG1whonB5PlReS6/pPHCFoEmFVOmQciO/R/9kObmVvK2ruBQWQ2qKI
DUSFDLxbfWlPd9Eb4BjDvMvP8TzWV6CBGhoWXP/H3WBjGAobcdkBfpwrSqubpPjdqsTdhHqbSy7C
4s8ivh0A/Xilh9JCA07Cqnf11uKtSAmgyczeMa8Y1jj2iExayKKV+HMaEkb7Z2XkIE/Nl6yg2ZDK
vWjGPWEpzxtMDnuIJxvPrpqR8wEvHD45FGLtyDI4P4AbQ1iOdetex0MoEQy2L6Uf5FGK6MQnOMEF
eXsiJhTut60lhtFcQQumT7EIgCp6Hl0GAqA957VT8G4lH6cBfjYte4CAO0WYOX7bhoj5G+RD9pEj
AhKV/AR/BefyePZtzSA8n3fE9D9AJoYJJAEy8tXXA2ChI2hbBdUAOD1upZo8e9hs72WK5jYPnaJB
uZkVvfu4umP2XHe+BKOxMYQuMqza5/0vajPz82ZfxWQisOTJPpZ+c002vJORw1wSSpva92Ev3Yr9
W86+z8MX22iwdvRdAp2lLsDxtsEqavmCLdYnusZqZ2Yke/lL1ypHYUvodK7ZSCaNStceob0WyiaZ
Mpuq11N3WkftsmnSdXiQIRA+7a06E0JGcAMlyrgy0GqIrT3I8qll8VyxQsFOIPaHK1Pk5UGqJHUJ
kgFUBaqHhS4lRP7eLVM0lAcDpSNdVP6+ARysCsMmn82XfPpuPRDQhjAX14bsnaK28lVAFvu59571
TgtHQoWE9MWnz9GoWVkSb/aSEOlSTRa52aZzUPA2+r5woHzCcSLBgTAicqIK93gUb15FOnyPzoWY
3M5obnoLQAF0Tate4js+tSrQ5xiCzfngGSHRgwrJSzzx6mKskVCejSaNiQUPRnrza2bxWzEOZ9ew
YAz74TuKQIALLPQMKtptMl6R3HBw9cFqPizHhwMw0bVRfCmG6/tRVdowLPFFk/DzaGAXZX3ycO+2
bcNdH7oomgqXsUBAET16+9Y2H6O3i10KQf0Brhmg+Mq0FHaC6XvL5zOai4O3PshCeIj1r5sW5SwC
8/DGiApMKGRi3l2BItOIEO5sGfYYpJJ77bXsTuSbE/z07QbvtYTKzRP+XK+YTEE3xPWGMY8ZGums
39Q1QPKM/UqYu8xxafoBKXzsT3z9I8+9fhOAv04lHHheP/Q4EQtTdv1nzGHpfIVwAI1/fyYFs46H
6YbF1YCJ8Mg2a6f435M5xD8GEVY3VAQqEN3e6Z3VIKXkDZuvXs5Z5uG9Ju3Ct5fu7QsWFVGxdSqk
edKnQITywelNbn03Dk4TAvp+LqVuGNUoq2ZFa0O61KvHgwrIw/KRvstSznxAYPybtTLhZiyBb3O7
y8A+1YUhP8IQpQjGFb7SL18poQCJyXVgauq8KsHCbgcCEsr8EbuBJdVgzGYqW2ILtemqPEuLhFnE
E8mNoGZPqOI9iJUVHjSqOQw6QKoVGRgjMBqymGAqQX6XMZM5XD2GjcgW32zl/2cBnEYC8rJDub7v
Ivn51S83ceOi0QJ9HzyfmK1cjnIg9vNyCh0fFSrzHIdkEjZja24kNDAffknsOcamy2ALOv+0G61t
GAYj0JH6Q9DCkuYsbgMKpm7rzXBEGes3pMlOlsWx1eXTeepIeMnZu2YJ6nufVSLkgjp6Wzodj4HN
XLdw/oUdPBKaxTpxsQqt2tjuYe2du0S8TRtcnfcQM8bh5eDb2xID2VBNtgjh6VgYi/2Hi5Bk8Uq4
P5CjgDGBHTJ25sDeIbza7e81O2XKhfP43W+nwXclryFiDw3cJAiQTPLGX6R00oWgpjzn++7VhMZ0
pqnt1lZ+L1UI6pFd9Ouw1O96Yf62bzUwU3q8xAFTxGKKzJb/U7xeRnB+3i4zTuC0ndMuHI90ISHa
omZOCZdEjRXB9GOKxkrjZzrwmp/LMncTuE6Rd2ia0rIyGSq6Gp+ah6UpgDjMvWBTS1ma+74TV1DQ
dPE/9aEs0KsCPsummSU8PHoKdGUmXcHXt1bc6EX3080Q1S5bQXzENt3B03ecEXwO0TNCo2z7EmuE
+3f71K5BUHypKzSUrZGj+b2fBKItit/+DvZQThxSa+iwhb/kKpDptbtMBqy2mbFLHnpIHCXuAGQ5
NK7PMzFpXrwJn34IeACefe1vJzcCrVGo09wBbu5p0StCbGM82OhPlSraI8001+TihdF4swQVPYve
0J4mTLJbvWcDDaFc36HyZpA8f2S40rfEhre5sZQLC/5xLAh6RdtL+fWG9Gqqxgd2FukY2uAn4/aA
fJktSkM4wrdLjDYEcpV4GhlgadYT78kKuchnwEYrvDWEWTArHD6IgqfAZNcIUAOhjqI3TnMfWbEE
UJQnJrZxucF+GGAYLrYcGC3GlNc7cTXIgT3PawN095UKZst/0NvG4jOU3oH3ao1KjY75nKe0WYIa
jWXU82KZ4/ZtXKQoOZ/6c7uGCquV0YphEcyypMHTyMKlWf+PAYdUIyL/uHKxnyCOXXggy+uDjMwr
fCxy+voJI/AHGuK7Df2qz/edqBsErkPJcst1IjXG1rKVjDbHiOEmRDT+49lALCth9f6vNdXVkgYT
SZpCW6E9yfDbz7Z37IcYs+JIp1q6w7twTqTJ2tBC7wCN7Y1pIN26Cf17aM568LZAgfvwY3xCRLIP
9vAHTK6bLJhmp10Ewsi76bknEdp6iaiwVGSMK9AquTe36H6sEqVzRcu0DNdsgD7Wnspj+iX7G1JX
4LsFIrXaWF1R7scterEXsEL4wnw9JSAaSlSG7rV1Szibb9Lbp2P+wLoMGIMhKBsVb2CAOEd6XfP1
3KbvtK4kIffDWIpChpaRqlyRiz3f2SVRYsXQf1AvQ1X/TcL0xgMe2ewXXIW5VgJZRuqNCP5lFLXh
k/Wgx2H10nUBa8idp8hXqVPuFIdfMv06dlc4PBZvIZl+itRoyu1JcFfUwWVEN/ilWkzNQKaOvGUu
EUQiTLQTcUK1xJiNd6w01bZg88ANGEp/R2TEltOePQ7JTOa1GtG8RK88TiD0vAZH+drSh0n02DFG
xgBl2Pvf7MM/K/RF3oiLSOMRalSAmVpOO51PWbzyY2Ri1z9gxvyUF7GhkPQPzGKR7rHBThiRxj8n
r65T6xXoMKT82UnzBnYNpC3X6LfduuyPtciSlwWPxNOOz4ciSKnlyhzvX3Z441s5t6xMndWbemU8
axzuur/91iNSxlr3bDqln6JZucdV8EhKRzSXJYw+QyXFXf9U5mpkxgsLyn93ufMYCQSa4WKAL0/m
WF1OQFnlSKMgvbR4X4WWr28oPdcR62NuyfuBTBeKttNbWxswThK9ko9U1/scSbYJrgZ77Wg/vqv5
xNh4ojTm3GiGQOsKykWGZ0pt9CXZO+7qD5Z+fY53S9u6zJTjBGqy3OVeOjfIqwNG8EcmAvPnK6sL
ZV1TRrl06U6AiaUdlhNfW2KJ0Z0kh1ZUHe0rrfW9cO41KJvjB92sSqAQn5g0+amCrZYzpZlhbAu2
YrIHIe1xoU6jV4gWVNXY6dflup9P+If0/Sy7+A8dgY+Pe3gVNGUmQEMYSTVOsCehKmR3bu4MGPQX
X4fPx8UxEkVpYo9bUpCFgKiPh24pOAeGg44ibeWWbhbb+WUf2hFDl5ZhWdfxMeE6wMzbl+vYhUE1
6HYosD6pPyPw7RH0ygWTuNyatAtO/JcQ2IGbljEnLs3gqPopJS+qhYnvFkGAqzMHfZOlYoBx7kN/
kIWf53drdX5ErJuMpkeKqaxpxxyxcHxEsD7E4SkljpSLzANp+EZy90DaUOBztP0qW74vOkgkHGZ8
xictiMuNkW+P1QyrYfePx6Xaot/w828tVFw8dQmBY2rl3DhgxJ6I/x4AlLOX0uIEe3UkBV5IXU71
hEgq+Ieih/egRIqVmEIugYACM7Ft1bGV7XIIuran//Cm550GCyIgYhOTSqZ5XqJVjdTNgwpeydf7
neSla44h1Xhmb0hrzxKJH+0h8jSgMd/II8K0jRdm395j6u9mOxrWeyK6M7XYWzFDpiukN+jTNOHU
RxQbOo7BBh3awBw67CgpEPVvvcsfN3Z4GSSrhF/Kh36Y0MAYE5PewDJMHexA4Zqw4nDh7jzqhHJt
vSVrNvl2+QCAwYqCo7F1H8Ud0legUWYLi70vDT7vGc2fs/lzNUlZGX1jnBU6/nlXSeJDDVPm8G/Y
C9mkQlUUuKlkaTZj3/4tTwlAUkzQdfVoALq+g8IokrEn/RqqM4SvBd8BS2xgBJejptwrMwiI5UjW
ThoQqKxFL7X+kYqUcLPTblFyq48vEu/geD0GDOYsSRHfzFosm23sCBEUKQ4/OaVeK7QJHEaoIvK2
/hDsSUTC/7i/k1f3jf1gdNWWrqfg/Sg8JVWuYF4kNpNqGjVveunuJesPWMaP3RJGkcrBgICNSd82
zScXllJUyhWzmHi+WNEkRJiDWeK7ubu/pVy1rM10AE7IBFkhYWY1CiJj95N7JBWhNlWDyyPxSvNG
MpJF84WjTVp/q4W5ULPBDYcitv5hyFf9D6Ip9IYBbcp2ypmIMpaA3dhs2xhAEA5CCVQDqIHh7yE8
vtKdHvfap/45zJD/tjWvNqypkNqhmNcCAPaO94Tt0Mf4axeJwAinUi3LZ17eaVjEnrdRnWV4CBme
P8ddPhPlJUw3KBuCbWsGtshldzvmriP2MUg/xzi5Xn7yfnU5pWhO7zvsrovtCst+7zX+DfFdti5s
f/6v08xYV63zUk6qDCyhbb471PoS837pS4UW6s27J0BvNRtQu221okr3aFn0mN05LSzUZmZrvrFb
/HOERpSHCRhruDt5JORRdmIAgDh3bXKvpZk1K8GqO+LBy5tnh9XSJedgPdIwpzoLlGRWIFUuARrg
thTfrwlKvoTNywHA94hvwOGWuDBuZw5v0IAWrbFulO9S599SrcGhcACUyDvfvgyAa20Zf3Tsul0e
dBmKF1GVH59ncKNE9Rzl4FXCIdixV2klhzopewxk7blOyQg6ijWak1ySUnPeK7HTL5sYdIKUpA0a
oDSU2xB1RJ/SXYIuNl6YmvBrjaBj/u8fH+mU+uuI5N8so4UFcSgK/G5wkrR76tXdl3r78pnX3HdT
8BoXAxcx/7+ZveD8chtWnSvSArNawHstIQCL9auXKUnuEMo7TMx1I9uo/WneAVOtpHWP2tHEsUSb
JvS3IfWww8x6lyU2ocItf3Cqa2mszpRMeHDJWq3yMws3jPOHwlB5bXr3fwDJr4V1fqNvkhS6BOHD
7QAqtaXz3hMfsx4eNSlPYLkpL2tZkwx7+nckTKkLcXcjxJBwZrJChzy/yEt4dEGANixGrFpI3wgw
yQp5+Y/U8wc5LHY43/jzfs8RE/iotGZBzM2/OXQaOMUu1QTfpn9tO4yOn6sE6Hws/C/H87NGiBxY
XWDN4QZ74KDDOEjuefRLzeJqw6VRuhoIaAVtwTFrtl8FFv2i9QLWOlt4+98/Uj7yLfOLZSThP1eA
O8wnh6IEkbRlZrgR/3zT7d7f3TM6D17LVrcZasDsblIcuRiDSvIwFCb810ZgRsWGlLxVDTyYOUy/
1sha+MBes4z51DORlk43Q/b7TukwTYuBRzP7ABL6KOBBAXBqddnkVJjFpYAVlqqmjkplDWHOsxeP
xdbvLCccmN3bQXDMQkfMfs4qGapE3GdiiLuED3dB0pUOhN6tY/nocupH7POk9UhG/RqSPMO8XUpx
yJtaIOsL2a9WL2sRpDMA+3LIWo+VQZcf224Fw+LELTjUPJrUFUw/cbb8wx8SoxnkUrrc0aIFFlfS
+NwNWq33RqG4JDEobz6R7ShqXVg9dWtAx2g/0G/d5T76uDxLT3HkoJZ3va++fUnCcnIlkYAoS5Z9
oWvYOoJJlPRezTAxmD+D46oDoN1dhxnTleFVU55pdKBXKWw9mt8ShTPxs3qWfWmoZdX5C3JMzmg3
AC59S3OKh6WtZ85DUGIMsHWRqO8vvYdfpMCPlkP3fUku7V3ZJQOQOcXjgbk5SvuQFj+flku77ADR
EnRQOH06kR2sQ+AJWRLVDv/pfXMJUJP5m9UalMkX2vdl3Nw+AuUfcoJhMshM02Nc2OF4XD3qiZLc
15M4jcwFCSXIAOg8I86LFxb0EbXXeF6ZSPukhPo31WnpM4WIp+f98Sx2gykcx+P0UkM1748gMUUV
r/Ac2/5W7SpbgXctwjswcrj4SK6SDtsCEzQjnByPDk2VAx8FGqBDdKenvPDILPcxS8Zj1E8CYNp8
7bed5bK9Gpv1N30MOmyzLIiJkuuUDQNVTaffRdBzBiC6aG28M0Op1yij4kmzM8aQNIECD7hLbN65
q6b6fwhVNm2Owf4vF8SBOdVYVa1UeIkgSNdg1bcF5fNXQg64mOIMGrR+hVPab1k36uzIBGTdy70o
F5RYqm0FlnBVuZTP2wMREX0sideeHxm4yba09tm+UTqWTnHEudaMrpK1cPZMoNUOwRCPzbOaHy6M
c1154zVBTl5SI1+RAamrf6KYfNEq5+Hxa85UD1A5v5TuztQMh+tRaoQ1nPOBGB7StMESooCpUF1G
p2HpeTOG+pGzj6mNk1ujMPjqNgPQZquUMWT3hrGpcyGTRbji1deN8tGrtQRFvVPfkSQX70hCLOGX
gfNGBjuDGmw5J9S8ZqpTZw9/78FG69VRDXCSux0i/sX80aKeVgi3l4lcFe82shKFUW5HRlax0+tV
JJbC3eYucLtDqzFhM8sjvoMpTht4g+Vb4AuqxIv7NXT0dhhzXf7SRlpx8yB/gbGRAlv8MhEnmQgL
1K3sk3kVas3BUFsxb1VzsWOgQbqI2XfBDwKFqlOaRgoIONBUvof/xK8V1XxjgunBgzTvdihD6PJh
uHaV+haPiW40jzXB2ujJ2LUJ9XJGwxPnoXJbKeIixsMnLvFOAzJZFeIK+tjas3eZ/tXpz5bQ49w4
lHSat4W88/jgsp4snZszVjAQp0gnqg8IXWa/AEa+aHLvxbKSrRfqyBO2RQDXsc12uTNo8ZeCPuUj
9WqjJCGapAsaZU1URaZBgewWvO5JeWI+oxkIUQcL1KhFmApB1Bvi+b0hpBcaiTjoKpjAUAvoCSWJ
dbClO9Orh1IDZZme98eDCpI4qNHdxb9xy1Y5hAl70jiIxdD2H6DjGtzdHlgVtF1fgTrv8fISPB2E
sn40GaHbyMkLo4tgd2D3gMZ2ods1l/+ZGtTiBCxjPv1uTcUDoPYTbgQAgWCgVSBjKPmUkVyrdg8S
vCY1vdEzcW0YOcxZ9R2WMKIMqwUnR39pP6ncWipZMS3Zk/K/Oiyo2pzdgDCiNKvWDh94RN0X4rM6
ZeF64E7q/39J6krpIjXpBGfGo9gLPRJBJnKyCTKSLTPNIAX19RkEODqOFGGRS0VjyWAkulfaf6w6
aa6S7CeCnhzFeHZgjeKSxy+ItXtU9uPwSPi30fZFs16plcCVo5kOivcs2JCIMgMqjTzFoCYyvJcu
rb8HDn5sdU2wpC8iZLqfk3bjFaFDWv/1cKOaEPIF1zNwMU+d8D429cmEotvwARMPaf2oRvgWzsHN
SyVLI0UyOUsdlsf2x+v0fOVXxxcD/nRkacQPiUQXN8fDUywpfznLO1mQcIFImjDESR0e3x+j/r0E
unXUNf9b2LbYt76JvWSNecJtgqRAITsBTR4U4dcUWVs1ZI/hwyeUcppF8u0A5rT6IHTVd/L8r9Wi
4wdApvjqDDcwrzKONOH1zwnHvIVQPGwMKx037hUhZUgAeva/SbKx37iuxS6nYfn1evkN4XAK0Kmo
IDpk6l9/s/ynbQ89ChVMV7NjBsehZEiWr5gPS/NfYPaC7alPikMH4/wCw3asppHqB2XPoC1KMqC1
sf2dXdmNJXWbMrKowUTSe9QIRMKCw9OsiXg+tnuBIwM5I5nTXc0SF6nUm9lxF0oRU8h0fzr3Dwff
RjnJ75E6JcoTLNDvqXAAdGQfitd0I4gRjCrnLZmApoGAA7BtbspeAUgEHHv1RBCcw2TkdRjtdmUT
7vQxfWiuEdpaGdOOJzjhO4gCnQqwS1tdMxsC75oSRJTsw3+gyN5vCEiPfBxGoIstCmA+1j5ROJ6L
F+xdP7s3M124CIpufQpMU2tUVMALydRO+BmXjd8TgBOA/6RpIM+twIHdS9K3gHWnFdY5CY1CEKTg
efLjkvR3MHg4xtqmhpAkj2gaplZghmEiruQJGDdJ09nwGLe/OA9S/vHPmtQ4SEDQMMXKO/4H5apR
K06kRfvPy6InuCeSSXjNYR0cM8JZ2WBvBzqitNRoek3yPdST4tqI5SR9SR3+nXvTfztCJw/nVeXt
fAB6da6PdovIkISZkIH1eJA9p0W0dbob+YpOlVyDEcWLWQMh8jJm0nzLGAzktaVol2tY1CBBeHnE
fVDolF4/cBNarR1SMfraTeDObyyHD1JGSYFeBHIzgNyRd0nX/3UImU72C+L4WrYoNKqVb+9x80aA
VCLX/wZ7ow5grGKm9k4/ZYC7FzBIEGG984Fo1GA6JVylCi5TD2jrUTNFJZwRlpQraPv55/IZaWVr
WnhqZSUddpfxFGTIUEyCfrYEnuGIamKJ+A0VvA3cxSJTmqPf/e9cXArejGkjORQreLBmEppmbLZa
4NpXrHI1vryZ2btIoIJnO4Tmyu0NNkPlxV/aYDjEbtQsgrOoGIODZfoZ0XfXdRDK34dFKoVCEijY
8Xr9ZFHA1A3K3qD9YfFpWDiRDH8uWkVzAr3S77hz6/WppmsS1wumyCZnrfQt9ROjVpVu6gGXnr7z
OvmRJPW5WppO0YnO1IeND4OY3fdTdkYBG+1cuQ/8RKidFnJIsDqibxGQAnROzgZfyJVyK9dBpH7c
GYDuhOHhqeRXZjlpwSl1CNzZ3z6ZRdR9ELKYm3bgLN44aRhoKbEkMhTXSJNk8yMAshl5eAAwPKJR
5n0Lg/ap2oBt+folPWpz3lvAVJU1sNi7n1EMq+LLE2k8THQiYpCW52HmZTXegOsMLtkJD0kRliKi
RYF6DtpggJhIb5oXwx4PgEhxc1VTvXCwdyXg3apE8doBc4eMQUELRNZx7cjXw4tF8FYEBXHQi2+5
/oKt/hk5Q3TqE3flTVfH4j4n92E2hjR1951TwABZKuNQDGJdWdJex0X6kBTfc1iUEyaGH21nDEMX
aHeZJJdiQcjNP+olx9pgun2zkuCaOGHkk97z5Ax65WmSrcHuRUpTTAsAh0HmsGLHDyskic/0BP28
bi3pkTcTYoRTzsdMZhS/MvQl5WlV5K4HBJI3WUdt0HQWcqYbmd563iL0F7T5cHFnFMAOxwgowcRZ
qrkXJ4Jh6iIpk9KnWffyyjWLU0NTXJUrcupIUb9RG/2eCPvFM0JL11vI80DVtpAqKnXyd9e6eyAw
3Aw4LjilcZkAeFOkQIU9L08SsLK4HjaGfy8dHcgxLPac1ocKFHyCJWAcvP0pscQ39of252bIwPKU
56L5AG9vez9fWtbUW0QjCMhTsqXXaOCWfVBq5oAZvfe7MH75WiEh+hq/rg80o17CZrSDfbTjx8IW
2XdXox8DRx38ZagEDlFU2Xb6jyLX8xqNsp7tKqhu927Mip9p63J0WFflg4LuhXldNr0+CbFFyfJe
qDOHAaaybBxw+m/d8MbgE4bjtHo+ePbSbFkWQmw+ClkVwBtQzDmhCC5yG23UGzWWmySppMhQ7rkl
DOPbU6vtCgAClkz66AnHxrWl3ZikOnb4HYVR8pYz4TGLoztf5FVs7LWn/ubF0A8Bow10i8/dUXS1
m8upNTAe1P2l8SsHgJ6JJZxTXn18ZyOne1MYD+h/fGGyBl76oxk3EQ/HE+7z9oI0dQfvyfVbBMC0
7TPbNl4QtnSo5N+s2iTShoSa4e8YV1/2JYjXjR2w0nXwA5BIUKuBiaf25Xs6q9JZYPnHi7w/pBNE
TMnd95tEB3eiKL/kN02CUuW3SEPI/gYu5RJ/8f5NLgR9FWdZBkYP42hKs3sn4nOC+x+kjCI0vyVV
jHuEbRkXyA/9ap+Kf6wSHyAVUJ/g6snYirDLRTNqE58XQSQ2klmMB3B5ltRavb7Bmw/EMLcYdnaa
y0v5OhEbQ4cjQkkPtJDg1d8VQW7+gzbCLIzycfUbEa3KBY9r7LzVUO3QA2tw30vTlk7mVwLR1S0K
Tyvvx3uAb9+J891jGv1gojTBER9tWREZyDa9YMlvGcAt4uAH2iZSfzu3OyxP+cIz79qY+oDZmk4F
cA8L7Tzzv9W8+TJeACJn647cZxtKBYgTUbXKWG/cpOikpj6jOX3/Qfs5VoA+Pm+bkk/3rkf6Fjyc
j7ECjMclV1m45WQXh8fvjH7xPJHu3Rc7svSq2Vrq8r2jqnMB1y4CsrHzrx7gtG7zBzyiBKQcC59t
cpZ9CptQxQ2UhPsDbJ/lpxuIKKViAOOxRDtFjGJvJRvqcwVrJT5Rjrp4PyNQk5O2Ici7AOL5U6sR
ONfnmPfkEm9iDIcSSHQEJl7NjAOenPc21OwfDfL94zSMSbXhXaFxg7ZT8/4neskKAZheSml77gBj
wtDYeZR0K8/wM7Ix+hvnWLvgONsiEKmKNPILgWhW7fwaztaBrDZGvwVEseADqTd+2uxMMtNxG5nm
9KNTZn8Z4h91HhPbZDygNH3o4dFmtgXwm1LSkvR+I9K0SFR/A7sjG5vi9CGnVMUUq3qcayF+/yZ9
4l5DDPnxWYstcCJPfCrBffyN0eXEqV5niNyrpWfAzI2M/Ke2uwA6Tf/zOoP9SmCud80TqkDONoW5
glomj/iwt8vsJfBJOlFzB8ZG+NIAH5kT5rQv7pC46RcFiM2TfKmJlmG+XHN7+ZdoMRyHTvPGruUo
ZPyVYF19bubp9TMLE8Kyg4gCZ5ODE3tsuUVG0mTd6tDrckeXtSu3Hu6QGAlWi0iIs8Vnwm+s+BQ3
q8kVT8v8lplpe3h3cDWApC7sjYKJQ9YTW4pm2fCMPi2N8GEj9SY5vjPK3jDIjr/YPiY2QTfmSerF
8qCjm8mpjDuBGYZ9tbbxy5mbYtsyO/taxck7MmqBlwnbVM9y5PXg7/83d27x3OgW6GffL7/kdT4Q
yHD15sRG9bt4AWtxFpZuF05eRuN0F+bUFO3y+xRRHLfWva5JC8R9Gk8mLQ4I0i76x7/xkHnW3Fgd
C1H/NGQea/Vp0uA0EN5h+8RWQLkkKnrIgXpiv7SENJPRW5lQ+ZGW9u3Y1PJ3jsL15EtIWUInGsb3
l1Gkhqxfo2r76nGmSSfFn8OWqXIHZFEE44JvhDYQ9UJWyBVkG97DJMBHxyX7RB3+s4qcWConTtiD
hfD6po5ik2NWj5Kbvh670OfUIyBoDfl0wtDsj8dGiWintN387RHH0IzjiD5BbDiqiLnpBLeFyP7Q
U2nBSWb/yeAusX1UTBpwUcG6nUKm+s/cXcb8tcQnI4xcI45OXCHOl6rsE6HKOPKkIh8S9DZdPkEa
5p59qP3jyxrBTps/mNt+n2SnCI3arDuHs5thDoJWTUO9f6tMADIs+WbQfgqbEdntJxoyVBoU54ha
C5Jt+Zy3QwUE24T+MwTA5LtVXYl38BRpiPuMXrZ3Wd0C249ZsDIUX1Iy1rv93lHTz4PQUWrUvRFE
D6ssWsNraJLgT9r+VOWSWKG2KVFHszQe8Ms00txDDXDOYWf+oxk2yILagd3lIh5c49LiBqDIlOeL
eP80ylO73O4BG4/bzPiZZxi5rtb2C4Vet3kaC1IDIil/d3KoZt8/DTcJ0uUDC1az/aiykPQg1l/l
5q+d9r0DXz530Hp7NXMXxlcirw3aSAYW0IUC4tsW+cos2BXuwNbSEl1XZ2KdhLiC5pyRtBKcYJWK
zepp0f/CWPws7q8j8ZyggcnxZB7JDA2fHh+bllv7bEFH/XC5YbEGwhKeLutt2NCD4szANuaIzq0a
74F1QKxV4vcGC50IZeAHL2+tb1cusnWQVJvDhh/kifk9PmFywi4xXTB2jzqzCl+mupy/jgCHxJZz
/ciNCt8l9CpigJPv2LaUHPz9WcP9glJl2lIGMP2YhTLm34SluelmsYp+dI2GpO8E+wldaqCKzNDz
acGFuzZfZDuLgEfyEL27aCtlFJEQ7MVVhdvoVUR+ZVkTlGqTmwBMvKtNGz0jtc5t4RsCtWoIslK0
DSQrlxOMOfcry5EHSO1aEI2Y17x/4+JNCT5yYvS6qcXvPEEWdtXTWiMyEk7iWrbA9QpoCrqOYSJb
ZoISwTkgjt/kfyOwlz+w0rQwvsbkMKDHTrgEAdXS0JT3vhwbUESWOXU3/+s18ODHIwwlFfL1YVL6
CMF1Bcm5lVj6e11234EmrMtK/bpC+P2UxV0k3UzB5FtvhIbf+0yd4h8GHujIop2wSUG8NEaocQaa
MxQgLFBRxr4MJI3NZFAg13A3CffXJFM395bVIMVWBUWH25c3FXqtqvCLuFAqPwFGn6A9k4YIibg4
m33Y0fF8soqyE/foTqaO3Q3krl6eErZLCXX9DEFpkifGkB3AbWvO32ChtTfi2EehgaehmqtzrW/m
XszKB9UO5ZAs+/L+LctDKFLfkW9EI5yxqL4gh+1ml01Ghk+N/tPht/VwPpCrxdIQWeewoMjnWt+Y
xxbnTpG9wQtfT2xIMQET653B8NGJv0QmkKbYGH5DaRjbN+HzGrpzv1B1mlU9PMpCOEfbZ4rE14Fq
L/I4vieAlR8lxsHNV37NrZwaKjXKmIo5iEcF37jUZT4uEUZfi2cQev9tF2WYwQnp/nZ1A9GBM9UL
jRoa0wRHC6s3En5dO8LKydo350RWR4DrDoNnOwtvhA6UGch4L0b2TsSwzfX0I4roYAyM1fJydiE/
pckQwPJqjYUcoTCvB7B2uw6G45eEzEDdgpICzN46P2EkOM8vgsJFBP8hNsXyGJrcp9e5nR0n1aYG
OFRQHXmScaIm4SG3cN6ZV6SJspF0TM6bbAfEXgWYbMWXd+/GnX8zW8ar4YNOzXaCn65hnpe+ffse
pC9hszOGyksWXlI+c3YXbf5IZxVCKqKUFBfOt93bN8/rXPl5VVl9Nat0WSe81s0sB2XPYIzDG/JO
C1amlghUsVaGLqZ/lGC47sJ7FQvUPYk4w3mg59yUAo/PZgRe8luZHqij2C6fj5d/NZwSaB7vX0rb
lr0ioEqGpsQYeUackIFndxxscoyPUdw2hxWjjTbyZmFzt+NTuwEzhVNXgQXNSDp9MGs6hVVs27/7
FXn0qikdHMDe85I2FaMRAOsfuzuDC9UcS95bSnf3pbwDqYrZnV5QcYYE8jw4CfIbcOOHVDkF6Y0Y
FrnPfy2lEbwxKvZHkup1EP6LhcrhiDzWj+IW+g7UZ7Myupy7ElFtvaJmNGyHdtpjxF44nkp1f1Sq
bpWd2C7e4xL7u2/2x3GEbi6gqRVg/ipQJeru5R6xnnERm9YJvHCzlsI5uf95IxwonW7J1o9aJ/oH
NxYP37a2l82LdCrWhQsmbU/xXfy/InhUsNS4YoTVzPVvtUSeXD+HklSZPqLN+Z1uyLUj8YHZ2mT+
juG5d68/pGCnYPy1tp8ZsVBn1ixN2zbxkv4Wz5g/hNU99rNhZANSLVCcqIeAOkQMZUiHbqSbgj5T
PPhHpN16wE3OnFUn9biNyFjKH42ftlXhLEPWNP5Z3y9YhTR5wdZiojl3khqxH0oEvDiSLxZGry2O
37ELfcvB3bg6TKOpXw98vr6PZc9+EfCEg6LR8hPyLxMBy1Dogdnh5Mucb/Yukl1C/6714yvqy4Yl
IIL+gVeVk8V/xMkJuJgyqZ/XTKSOxMqJukRJm8R1imWl+1MH5zSj2WXkUZcvqU7JzLz1U69/uMa0
N9Ybc8CFQx7y6EFZzmqWSCBGD7yQJ+zO6Ui4x2BwrHbmWVa4ksnczUf/GL/oeLDYoYAes40MZf3C
mb772htr+hH+lOhz2m2I3JJTQYDUesX07pSA8RznUYn/a93N5QDuaPWYjFNBFc+jAd6wvhI8HG5H
LymAS0sFhin877wKpp27xW/epxuNbjT+XHvFkt30GvzhCEeXtP+Ci0Lg22AWCgnpbe832KOjK7aW
Z+dtUbiL4JRpdPTjaulLYsfMW0SF1N2jwglB2iSWZSyCiLx+UdCdxiPVS6pJWpDxXH3B/DkO4bcr
g+XzY/Sh08vfgi98PLW06IXUaVy9fSkBZIkh+F9z96TFIe4IVrYVetHPrCux64uIM1yIsFpl3REl
ipmbT0p5dfF+xoKrAMzuF3Pig4DHXCWzzM6ukdivGs4AsDTxmKuM6BTnufpFZxYgmWZD/rK5uXX/
fWr3qe3koMi5KFTSvo6yRGiQpLNqKrnz2h8uBACITRvmiBoxoyxb8TpLMvfD0sltFXOlwvp5Ffhw
dDTWlDjJpe9jVWQVOtdQ9LoCRAhGf5tJyNnt6enOGVn+w/cuyx2nHcX2lCiYrrbTB4cy6kiTKUpP
Jo+llvdPSywJaWAHV4mDwuJH5AHlSqCufhL84tgq3t8fAXbJgnmsdTyIVLnII3C1IFab0cwlT85+
o99907j+cBfVaG7NMPhnndmy93LJUt8WccPJO56ti83KsEVudqPdeT+Vp5iAKXu0Q3dQNN6aSA0s
sWtNGv37sLNF79pKB71fq5Gjqj9MduDuKp/cV4wL92hy1UfTGQ0MQY0RMWvFXbgkImgsIIdZP99H
iukRveF22wOXi2G1jATzHuZRXfOBBy1QH0a8REQVr8IDkEMDCjkVl8sdNJ1ktE8O7h/m/yFerrgE
yFnBMjaxZyNNzHyPOQCJsGmebMxuKf6UnBZtU4qpPsJdvEZXwG7Hyd5/HwYlkk99Z1iPvkdHlws4
mMaxBVTDRYPQGaXdryoemflfqXbRUlP5UC8O65UQC1Jipfr2Fihu6yZvhWQd2kVbXLN16WqgTvGo
jEKO/ywlHc3PFPTQeQfEU1+dD/xrqnnwfB8UqXxtyeOCNo1ajs0BsHjQ+uMkl1x8Cz51o4jkDB5C
dGutM9JMCzMWXiF2UF8ZxXJEDKQ4mKOyqCxDQsVFvGuAtRQeUiXH9X4q6tiwxJnTyFRKk+ibH8mg
e662zTrVutzVcSSs9lGvKM06BX2UQZW2fexNTf9MMMBKfW7g/l/kq2aWIC6gobMn0iUBnPKUIYpD
sk8xAolUtaIkW5Dx/LZI8/TROh+BpXXOScEC/hJU6jvsmOmFPlsGuTcgh3T34xYmdm3NiMLXCXjR
hFhtmFNQcR7bMlLUJXXrfik/GFwa0W87gNX6mLQb5JuLWdSYFIRBT4EU2rJEh7/Kc3XtviyfX+GF
dVJk7p3ft1s+O0Kq5sFENzDr1ZuaMCxYoDxYygQTGy0RSjASRbaC03P3uL0dkrJQn4YDFY978dCl
iXU7mPNIgB3hZJX1UTPGVxaiFpPUudF3mgMtccdC0/IIPipjQGYHMElI0MITNNYttXJbMmliMI+b
auVNLtNMmHO8Rvzd2lVMhXLbRPTX7dd/oYQ0n7VzuPfP+qxRs+a27WcB4qwmEDL7Sw4rPLHGgsHk
JL1WwM+KZF6QD3faSqTJ8qvEp3bohYAWqxpVhpud7U81+0A7HJx0HPsI3keSJwh+w5YqgpgwGBSs
9ePxu656F0M7jeLmgBbXttFOACSpTb+PrT4EtsWxXkzIXwvW8EACdkKYO4zSSXzw3eFEXlhV26uD
cPndq0H9wJ/56L9oo7F0O49I4cqrzvDi8mcIe42yGkiDBD6KEAsHeVwKI3pHOZo4kHxlaeQKwekG
x7x1+vGM26tHIRXZ9h1taM5uW6U9Pc1P9YRAN2BuQbPINMbOIqwNbHEWFkkXI99gmCNCdHwEjVey
UXvxvO0DLVRHBUjypZlEnqSmyvbIbot+j7bOAm3sJoHipq5B2zRQyGN/tyoI09ac4J38Ws6fP5Sx
RLAu8oQXQ9vUdDhu1BMqZRONOTMl3Yc/gITu16zCNItpSjbwHQ32mFwKdzCjZ0setTgNminUwjpX
n+/yhbPh7YazTisAqVv2R0QWD6ebD9Q47GLwfV6L6SyA6oYLA35/kTWE5B94Rqz403SU2VQIjUHE
KYQkuW9f+YN/14gkrSvMYqsp0Ce2QhOGHnEZNv52MZzpfdom+8xZ5I0cqrHd80uu3KuTAhmjkWi9
JmY1elo1UKWAPmOTUiy4zhVT27kKkqVEJvrpQl6zJ6OGXnbhwyo3iYFh606uzuUDjawZ+BoQN0D8
jbF9cuTKQAeHxnzFCAISoeVHTt/Nooj0LGcuy4723zxf84zJY8033lGd5qSkTSn+2BEMFHRF2MHI
+kI/49V1Suh7RKR2MwkZSjdhwtzmBU93dfB17IXwnE9V8wdjY39TbNwvHW165Gq1xBZgrFEnEJnr
00tngGDYTp7j4/v57rThHQDeG3XgU+cY7ZqmCnOB0VjKL2hML8/KCLVWbkL/Ag2vz9nzXuNkL4Bv
nVLJAldZhWnCFRO7nehiqRmsEV9pCfjF8wIVMt6OgsbGQZ0VD0PBXAB8exh5UpWcDsJIXUvHB+RX
NC2O0aSDxNaIRkV99xR8Z5fuLcQh/COQfL/RCGVjhDxq5QrWXVCRVgFdFtFBh+EZbk+xzzfzJLqc
ZueckMBvWd26Ghqj43V0Ow9ln/c4ikGlUrdXrzxG+QDjk9lLxVPAKqfJuXrtM7B0BSvzoVFi6sF+
rk9R6JDngX6o2QJOp0tUBZjRP/LfBbCVuUMcxHkNxQ9YY+qXSq/a9K3OlbhdW4V3tn7QL5WLQgza
2W0+SbjFo/CzRcsYBpbXCXF6GrHyEmiBff6OCOE+Vk44bdsyu4ovNH1s023xp+8hyHAV7i2nEw0p
dyjNX/89xTpCa0IIM8qV9AAxBGLJUTMnfOHLMwg4ykLeEQmjdNxfL+iZy7hhxtAxcA/OXHIGpG0T
qFJneoQLpE6/dPtqjW8m+egjWb3eugxDnxXuCQgFeykyFyaac4tDqjrORmUL/uFHIDIMCjqCCkCG
F7sHLJ3rn8pv57bXK8uOVzx1MQXmKuu0gZxh4G5nJhESJ39gnI5y3/U97k7Z+CWOOF8lfFbzUvbh
vLatHk74MezK03ayhuPHL6V5pG4wuwvHMMxcisvEBSZ4ARXde6pGw3kkfNYsTp732H/3GgRhNpsB
se7twQrAE4BMqT0xmtXE3nmSNlipGb3NMTP8t2nP3QEeTMex4Pf9bofDFfYOhfButGCDNyzIILa1
jxzsdiyPTPgwMg3R+rsV/11dU5zSToS0gEfAUhIWR5eWcNWdDURz8Cp2cYxfy1Jz+El2t73u5pjB
xdhdOFfbs0wOS6lkUXgL4psm2T4rxsVGcgitU+hvEMVnljxy2sRh/Gru9Tla4F7ThtrXy26bAthX
0/suUVpqO7kwe09wsXsk3dMUgz1A18B9bheWDjrY28aoJ+aB6l40LX+ELezG29KvMSNtqi49aUAf
gDTOGfcVPPAnLA1sT5SbJoCrcYkwRPSkJP6kTvubgvfk7X9o0smc/aeTNMP1QUcuQUlPcqlnDXVq
GoZ6I4u06K/U1Mq25SQswW+iVJOy1nP9jkQN8BdlF9WV0UjooC4ZZn5iYhYhcS0RCmTozuJ1cDp3
vp/XB0cwS3F1jNQOLQtcxJJ+4MbzebM5NKL6DAG70/aNhadu54zP8129pYXhAcg/DgwycUnzutPf
XROS6QS4fYxeaAUCydNgLdTNAbMC3cJTf7tinMclM/EvTwSGTk3glzue+/cQrTQHq7MStmTW11xW
avLJsokAyy5zK0VRQkxoY9PRPONB9jKFqVnFo8Glh6hVefaS5HratGgrlROpKWK6FxmAIebkJVDJ
j+RCloCY9KQv1Ifz61Q0M9tAECl6EW3sn4Gtv4am7aEu7rvF7qdzWUBj/XHVyGbCSrHUtnH2SNw3
GlIdJr/Tmry5UjYi+I8M/iQq+MaJhvaA5C1D1TsgpuRxLMpf5wfx+blQdJWtaeCw6ne0LbuxHHwG
N15d0t6tJAyyt7NXjsET64DzNcq4HoTg/u/BaIXZPWXgGG4Ll255JJ9OYlB4Y7/n3t3Nt+wIchOt
BK+nma+JoFyi4cbxatJK5KrHN22lTs8xXPAj9/1DzyXnLz4lV8lgXKKy0rQhllu6esNu/+tQOcNu
Gd2AcWicO/RCHinX4a5udPAXmmGlPOykIfe0nr4/2SuuBNCyR+50bW2NxhOWYw+E1+8KBcSbXB1p
cIIGbZoGWmWYs2Y9ikW3e5LjJUnyBSiamElQ8s/+gh1xNQmkpaXy43TsHyqCnxjZnor9PyMOcMdY
E2IXGijh3fOD0F3NNPtaH5x3nQ4dvHwFpV8wqw0AeihF/QehGU+RvcLuAA3/hIXGCoaUFIaV8jtt
C5F8MeKZ5cl82JMLAWvrUTamdd2mNugGqkGwn7sEapOoefG9Ipxcefk/BPSMBK3smwdc3D1ut6mt
KkoKAryRmf0mrJrw40BFoCGPbi7A59mHwSHG5o2z/JbaMPaMYv5cezZpjbG4vYsAFiH4kW0ApJmB
SlyKjIw2QUWxnfQDuICH6wkA/jqVDFUtudH0/kRa5Wh01Fs7XK4tWC7EJviMLz8f55MhIEA489pN
5zcCrloEbHUPYAyeMVpRsAYww6NW0tILD0fhMyxWJhEmvYs4mrE3wHumPrZwb4Ct9r3W/T/BCS3i
YDhmJ+4oScM+5FZl+D/OZEqaMsyLeREuvd2HSKmEUzcIdGdksOWfOjN9m+Ez6mcPUaWo84aXEZS2
3WXFDB0ehIc5bHoG+omf+fd4yyEMqTM70Y4EFXX2pHZGc/Om7+4RfJCITWE7vz9Oy04AvnwaJxLd
GgKb+5twbXjd6pPlCNDuylatktB1Nx3cspJtr8c8rV+XL5ebvPp81Q+CFQVG5mCvRPitd5HKS2y6
lik9JpQp8KqJOEcU34gD0GLVpLo2cMFCzZcgxJZeCcv1B1uhMho760NH8OESy2Jrq45TpAjmiVd2
cyNZIxhz/QyOH+9oYKse/CX57YArJAAdPGk6TJ5/YfT6Wdg3rJYL1fiRknUyho8xKvcOzoWW2/Wj
dF9naY201odzJD3FklxX3q0xJ0AkI6HscVvQZPmBNvqC9usKkKGGVBROdkAQk3JSFGJXGmmBafc7
7sOVKiyxBKMNlDaymsuX3qxP6OEC5Jw9cGjug9Xb5hxyT6xf2LQLtAyqMTskJmZBHZIhDU7xa7VI
dFCCAw7EkRUVzzd48yPSxJDXiUbeMlbecJy93RHc6tZBK7W2VmY/GEQ6yDYmqeHPjCEf7eWaItQa
dt9nRLv14PsF2rJs5IIYADHtXUWekWpJApaffMCN/W3jGLb4GfhdfoOr/MSX2W4G9LaO0fYkspQ+
+thxvUD2xCTODrXKJPX9n0fdk1crL0uQ7UnM6LB1q3fw209MJIoCnAOJJvqQJbF07QpKXEcRPWIx
hqBlXbb/TQ4sMPRUa/0GMRFbayaA8q1cArwmIX2oskuMTuxTr0ECzlXsT+OvE8fHHPPm8bKkYoSV
dR2NBwBqckdlkOvUsmZXOV8q/czG9VhRX4yFlIKd0/NaZr88axdcxALBviVqj5sv6+qzmF7NSP3w
lB031BG7omBPULVAOGEKhOqjSK6VjsxJGEd/1eD+UHlMkhozFNW9tEmnEbSke/qlBR6KI53zki6T
MSPb+ugu8dW2ZGwAq1PUEVvsftKGHy7XF3VqwmgnSg06gAWC95eANz1U+BapVX8GZ+ms+NKB9LEI
+PR+CXT3SUNkqzcAePK4NJXR9nCsdEvefvew/TaMHRaeT8+XaGv1KIc4XCrDHG9XfUCtq58UsBZt
pm8QPwxu3fIHywNiULdSbEf7NCnn1Ez3VF+TzzBWpX3rrN5hZ9muKzGUQPBOvhC6YXsbr+qXomFQ
1/y2XGTpmvmx/+cMAF48kGb8M84x6I5zdEVXr2tM5E3+5byG8fxvlma5MS624vVCSeRhzHQLUJhg
KaqCCMaI0yXxMq/cy2CvhG39VWk5Z0T9Hxz/8xsijmdZVWeCVCkStV1EjEYMMKFvTtsbCaTsacCc
3KhUMMfbIN+cppF4v3AkKGt0arGprdMqyLuWeSWp2H/6ghCseVJIdRY6T+sBRPbbdTYuFqv6Isod
SYd8+5McG5JXoeRD4NdBBWT8bKo0WSKo9ujiNHw1IdPjvEah1gZyQH/Wh1+/R0v1bIUpEuaTUSfJ
AuJun91pIm/fgbwh/zQmRkXjYzFJl8YYNOoE507byVphccePTi4stG5Jfeh6ZkXFcZyvDGdBkkKP
mJBVDZx/v81fu6Uw67JSDf1HFc5b7901+BP2GKEBE+pOTUv8wNzwbEKZiUQOIk1z/n/PyWLeb3ES
tloTB/ztpeGDGTjJmkDX/wnl6ZuWy/93HlqnKc1p1uUfLFb27r0vs5FuhaXb+/YQYle1BdnJgCUQ
cezOpAB9hHVZcbP2r9uHzOKJzaGHfjRHjlxfG3YBa2S5Np0213388d4tUimz4EClLOP8eUa/1wL7
n++58FtA0Eo1GULIdlAzDhTA/caj+vOpycdgw3SCskWQxQ8zc4U81y2GE0PyFeNQeJ+mnN+eGcpw
LtohmD4RQnpGUttaMTVt7jm0iIzT5ef7bjK36XzrHSzQ3wdQw7TVgCgBsXVWJIYpN4Sqh8zPkuGc
9JWAZR2NXfaBrPsjgCDMd4iLxnj0Y7hubjKypVltDEXqitSpuFn/OAw9fPIZojBsDwVZHOwL5Rvf
Ioda9F1fAcH7RDCrTHFVwITKqAM03gqY/w5AR8GfDuGtIRKGLbrvSZKTAWyXXa21S8f0gCDeqd88
MwCi9dXx4uhO98fRjryHA4Bdc7/LNt1gbpIZnHW0MrYPZmbDfzfklMYIOmD031G06FuuWv7He4tc
NHIJdUUS4U2kvdYnl3wd2SE/Rzkqw3xGPT9RfWYa7/QAmgUBT5Eu3ikMxOGgMgao/gRUkXtyuSaq
2PZ1NwrcvoErfwN7YjkDmE7WZ1wO4019ryG9K9p9TWH5JTKDUoI15MaXOABeXi+Lau725W29UQFI
T7Djp1utD6LNz4luHklYRHMGAfDqZDan0d/lU1rtdV4tFp5k6cWuR+VZV+l6/ffSu7Ht+btjNbeI
GS+rdVEIEr+DfHAVwIIovuo9mXwyn9YfcFo9DJbjVofPuApEbr8xiDZYDpEXDbbLg9vHoT2r718U
Q0MJSV/i37iGu0cwe4m7hSajMwdWEEBMFN0wq+M957DXsTBNjU19dm+2fWQ/pLXq/y9mDQpCnhbL
YyRkfIzlidL0onCIxzk1k5AklgZgPjc++6cwv5VV1GILrByc5IXkLpOioUnKM0SD0fcS/5OnW11U
gwpFsABB1voHv/iPw7R6Y/i10KKRaARhZ9hTb/h7HKlShnaxD44/XUndZPxxMIlKpKK49XBmVrBE
VOjFLk7AtIJ9D23dLpYlg5ST/mlXB4kt8z6dBbqFc4n+EBM/nz5o4UQqLRwcR8lY+vueFNwcPiJW
1IwJov9DD8Y28Lmw2G5syjZzc2Et8Bg235Rue9tBfCyub15dEAP3s7tfH4dgoDdfnWgp+HbU8idt
Jw4O5Irg7ginc/RvGro+z+I/BydjUM+uCY02RBrNS31jpko4z65wEVVKpobfK9eY+KnCXB89wO4/
7syG6ttNCaKEe9ZR8VvoAKvvuu0QH6h/aTAIeRqbtuwlcKw65J0uxYid2yBj1pPb+qxLH0bpHcLG
PF8sNZSNWUgdxUR8Ds3jq02wYxLYom/24yiY2JBLaqQNqrlul3aJjQM+W/HHyzH0yFaP/IYjHnq1
tBuTWAa/xIa2vFS4TwvzoMEuYq5UXZ2TfBEKEjAh7r20RO9Y/8R3FPYOPXaRe8ML2RmPDRxa/FF9
G6/EgtevESuknsXu/zvWCmHdTYrDZMUwwMmpWRXGoHQtgvR5c+9SeFf3NuZ2rzH/8gIhHEtoKe+K
syOVIuMh7y70Y8nRsVfh/5k5YgA5b8GBGapPPJ9FxyDiRP3lJKOKb412BSyqcMeAU2+s7RwpFGNN
o5gC/+mq8T4R6FD0XYwEz1VfIcCeqQTk3nxBgXM5gXjwJpKkKmnI5V/tY6pcNOHSWWgbWPeDEdrk
TR+hyImwA/RKVxw3Ic1eDwZBJzzxNVwd1B5lbGdOERERW5TkaDFd/PH0pVUa/hQ0zFKSVBAgBDX9
7ASxUhQDCJ0VmuVNzVPbGFlcUZfNlHmFeDcX+tW1Dn1WWSQku2Iqwn1rfV6w03RO/DlkgSwW6kdL
U7bb+GAkepsCrVj2FQPGaGw8KWtFEtxeHNLhwV7WGVe5aCgBduGYr9CLBxs2xbTm8BbATGTwxJQ4
NMc7JSsyrvfiSKOs7pXIlOigvpcxqprmYRTBqHnnIu4teGbbTj8MYYYfBECmWUa8QFo0j7PCIiMl
zT2+5BGfdmL2+G8rbKyd9hqVZ/FEB7MIUy/riAlyYTLhaB3kzdn+gLyCMhBpU/vdDmd11GXyNEvQ
TpzLoimKA1NOJ6vU7OU6e3TDtgg3FPRwx+RuZOGKDRjGIilUMeudctJ9eBoNMvm1jMNDfuVtm47P
k1HJL7HsaOGdNpaJd25fT9cH3WUrMtpI07Mp1YIZDGVTaLQndhZWY4tWiuWFJVx8mMiQVI3+7zQt
8mwENQUB8vMFxAW50aULc9D6mc9qa/pjpOIpsEAxjk9kIJdNygHb8CrL78MDS+SwLiS7TKupYpbz
UgsXbG6CABpgO0WNGc3Zn6RvscXzguIlHlnCQB/xg1qJQ9lLz+vK064TCV+oHHiFRIhEjuWw2Dqd
i5Ex/PpEby4KRVNK/FAinSpT0veaSljAqKErf0YQXtI2tG+AuWQVOrdjyaGUBmPvQ6Q8kdkXzoPh
WOPCjiVS6L05Fkbs40lm9uci4ZvMlsOia9FrFdNM8DBDcc76N04vZxzs3+t6KewzDntpfPtFtIET
zmW4BctSEnQHRAXAydTKE6hObj3AMqhmW9PFiU30GcBbybFhZSPnZZTPXI+CNd0JW5o0GuTRyBFV
2IOpiWeuqJ3prNRyzjMedHGkHfcT0MNZPo9zg80Jpa7vbWdSoLsACog147M46e8PuHhrPmKOzCOX
71lb/ZpW9Oiqp7GibBmGBGLhhBi4eND/WgRLFrIOGAGGZcb2znji1o0S1T+VKQ1ox+y7vzRvV3sn
su4596nMfilE/PVsyQvHJDn8KaW8YyNrkx+NMK+lXWVCItkeytWaM5UpbVUXHDsdVBk7Rrk1gEJV
GJy1QM3ebK9wSJXvogxLOhltLwqYZlKBamfyKNmuZYxMX5otgyTLZx8ELb24zZJuzYCwwOzRMcCg
VI1WdSnK+K7QOkpFgLc7S4WOv90cs3eUa4G6/R7dT2FlfysntyZxhO6kYOCRwLrpmfvyNcWrgo28
euXZbN4h0EeV5ti09UtAdw54zZl0CuvDy2+fWhL8syNW1DC5MiJTcGFtUjMSgq/+wMjOsXZ5Lj39
xp19Jn+4tsFo9F52MevyPWxWPSfSSslm4i/QHwMu+Gyo3aVx+zVDXL2ptA27BcJN1W29fIWXfbBf
9uQTdOSszkNsaZZ2jl9USW4DBV3OZ/rtxzHucztMXG4t5jtVI091uqMaBMYsBswxAVoaI6RaLDAX
Ku6+Un3O7vhRW5pzlvXyDe5qfSZJQwd8EA8+XCPd6bgGPjTk8jnGyz0zZHRt0T0gyENAqDYj1o1I
QKMgpfh/kByI87X9es0H0ae3V9H4xmB8+uVTJMgaMpZ5EcJ4qtNgL1ietgQ1KmUbHTcjfnvqfOm1
GotdUwTS5lNZqJ8XATO4acmQkH2S3nJGkdcDl4X6QNA8ErU5d8jzZCw43NiMs6HFPgeQoPXiarXY
K9JDP+/jJtcl/ev1vedjjJs50k2JUqr9qeUbKnmeWvKQehm58BKmGfK/ebSXQgPkRRYMJvUAkEfu
yNYhK/WSA6xuDTJ0rkz4lm1TVoQs/GUCHS05fTN325WZ4vHU9wTOSFvripUoaO3yVaj4Jabu9djt
H4howwnX7hK8tAGl0KYw4QEJA7uSESEEJVuQWRSJ9VGKfQIavD+lAxnRaKK4BvGszFY5ZcQHpRkQ
wcOyRLFuaVo04HnGSXQCgrT0xATUt1GtpCMm5LfIvi4aLEqtPDp0GIrINSo9O8hfqkWXoWMuJlz/
7OJpzdGU8neA9f2WBKwWv1LzaeHkcd7EdYTag5/MP+W85UFggmVU08ylt3OqHyW6cJWVKwNH69OQ
fVydacYW1SxhEeC+zA0pxnnvEBvQg9r6JYQ1EZ6fi/GzEOolfmqZWtsLeSVqX3CBc37muJBCzuwr
cBhNl4aGdhbZxbt+G+3/GD5m2tsha9yznw3Z/v1J4OaJ1Fo5gj8s6JM8KCuJMmn7nmkdAqnsZZjU
NsqepRPqvuW2/gh3fR4+7KiJqiUqWiHen6ETM7xizuhbpX7bPmRP1EK+APkThRhklFhI0goFyVak
T3J3FbuXzBxGtaMm8wZTKpQgQ+gTLo4bET6Lz+zWgwFG2J+S5lTAmLRZS0ot18uOo+6hkat1IRQq
zQRYBydaXATNICbPzwt5hXbI97s8jYmbvKTLPQzmz7fUgpcQcN5PSSkgcANSWPmBvsE5fHRHKbO1
ZLz9DqsOrZwcrB+EJKNcjdv8L4Kfo6AVqrysb/DmrGSmY7hslATCxuz+s1wZObAu5Mun8nGybNHt
TqXjneKlqETKKJLIr1/nS5k8/rRVhf422jQElDzQR0bO/KFBN9u4U8nyhOW2qFPRAoOzTDX9euQq
xs4uJASbWGszVbL+zwJg312EgdDWEMfg4wM9GgaqdI8KLSUC609nR+Y1y+TLM6OX4qOyLI1x29yu
4onuPD82Hgzg02wnsysleWPdnPQ635RUgBXqswiiDs6BDB/jkoFgxF36OELgjxG8P75By86M3XcX
vRToSW+APq9QJ9P92PPNHM6J3pRPCWaAVsf+YJitCYPoIi7Dn5OSoSVylZt/NEKJ1XsCbV1HRhD2
DKyM+bAfWx5TpVf3dGrWhvSr1AkLik/47ZVRKPAJRJjCN4QwiDT32RP3Ft7wZqjt1jgsuw+4Wrki
gnnRwaf2U6HVvO2+Wo8tThELk7FJlgR1cif1yQqd43Np9v1pNJujcElxm3H/r4mCZktaTeggjWgq
/7o7vn+qbuK3MiDpD5U8CL3Ywvf5OKYJX8o15pHcVEMZAcCbaIZ875vNit+aNZzNJs07q+MNohS6
9gzLWxGSlrotCGXYOQGsyykVILFAtXUBPsVeUQHxYNOtrqsFhRxiklGAd9/xla+2tlZQF/iUsI3N
Q0M9UC690nGkxCh2NmuesmOdVYr6Od5/b7UbQ7ZgftXKcFzJ3UE0R3N+ueu4/zxjhF+Xwf1L82Ll
0m9JYdeemrIczBY3XVeQB6yaK1QbWgfmx023M4XYXEWLX5Sk22DmKPRDxloYaEVs2X6oi55gyMc8
+4g4hGSWbU0R2F+x0IGDK1LxlDrjLsUtDayx7wSqda/BvThSoB8xrj4jwNy3tunlIa9G9ronnFRg
Qe++1YBmdrhRGQbBk6RMAPugl6icBIXfTZrxyjS/Ws2kr2NBgj6GeeGokeZ77Es1axK1kC/Mmhtg
P4YLAouPFChUXZiWID77duLZpYEUDO3A5qc3TrBGK8dX2YG4jP58yu1ibZdtx030KbdlRDYuDRdP
rkO3vSEm0paV7MPMioMWJr0PdVRBxmsKT+J9mPQSmz2facv4FloEZAMD0jejynGb1t9rUJ2BUZ1/
Yh59VqaHSv4yqoHQwIvdoWnMDLFdQLmNy/UPLNprWgmoI195pBsogF/Ik3TFNeIUc3pC+/0Kg/X6
V6UEmY7L1tBzgKqHYq1t5vrjKhXrASlyjWwFAtnByUtnmNhPfjTogNHxHbo0Azrj2vpaobGJR3aL
hsBt9P1BlUKkgeYOV6q30ZGz131t9Q0+aA8TX8yQeVy4/FGzJikNMAaiGROT9okR/zq1bx1R3qIB
at8KQ59LdGF8HVy7KOmB1hUuvGrMc05M71kuMlubfU3Ic8DQLssrRUeyf7v+IPghT7zR5F+LjVOX
577AhDUCbBQMi+Ev8pnv3GOYCEff5Ay2hTFkbH6fb5rGFL3BQsSwx0ZJ6G+rT/Nr0Y43akTkOsOg
ppwFztTRw6/ri/6XrSrVmFbKWnMOuiaa8iNIf0U4qd5P+7AcFcAkrdN7uMz+6hWFvC1B6YtTi5O/
kMfR9ZDL1etYlUFEngwWR2LlJyivcbJrbQK9QKwgonhuLIuzv5gHYsOp9pOL0P0O+KR90EUw/rQb
brxXiqt6cUDWqYTzytQzo8wTNLbvUsH9Q77nLmSSDvRDqxBr2VK63j466R2woZCc4j0Qh/xb+U9j
IKZsiZZZoUiP0m69ZfwpkjG4HZLbA6CcxAbP0a/NAfZcjL3SWFpJPID7WLdtFW+CmAVD7KIoUI3F
b2vkoqazU0D41dePUUFBder0VWwb0zOmeCWvSRwb/UlReKz5XZbfRwp4oyKB+p9mCbMq/Kpq2+84
/KhDmVb/igcWa7dN8z1xaEbiHiVGoCQORxaJ/OxatednrOSgOaP0BOFyPwXTHJaLDYCpF9Fijp9m
Yb3EnU66t7R3iqDAe90cktjm0LI7Rdp0SACoxtSjByL6cjyDloWa21uJOWw3EbbiOjsdNSxJR8g4
c4nnjrnYRipRk+zmnWGmVU4Rz0iv6k8SQpE3lZXMZx/ItE8e70GHOQVyiHDEav1cSj2qD/t9bCQq
oZ/eWmvayART/hbHOT5RlKYFeUKsnfgTn6uX+hjXptxaWldDmxhxE4NvwfRELkyOAVZrbswC3qO/
FJDLWmelyjgy1YQfcOTvPGyiwmPEPnKrfLnhzHYFyu0Ghf773yNTbGJuIQkOsN3PUqZwbuj4GHWy
e98PBqqA59Ex1PWsd0T69aVs3C41HBAavOZzV6KdLU59ERlpIATwJ82xRcXh49EffpGE5vqVjwk1
WWh+BQPh0LARhuLypFuLljgtzlHZBEEyNJPGw33/0QqWzlh6t4n+Xg1N9uhBkNbAYOTRaUayyusJ
WarX6w61YW1LuXhSXo7+Yv+odNAijjVk8DhXS+Ww+I+Ja+sOuqTziI3yT+/Jy1JscpaIeN2WgU5v
Hil/iH5eUhxit1oD1JdH84VtXxhphHPK4is5k0bSxYlklFFhYW7nGtGYBg0U5FoDJTeE3A5GDUBo
xhA/47YpatNXabuokY/okYaspn213nISncz7EWQrguYM0nX3tYUUyQziZQNaMEde+xTBXLIOC9a4
vr2F1kPHZIK/QPw2CatwGkHpHFraP1wm526s6QC5ZsQAIW6GtPwPe/RZLhr/jObfAVhPOgFzVaL8
9OxREIlTEyuP10X56uWKllnzVAhbEWV9N3Xedu6bPrcjsz+8zr566G6x7Ej3BmdTSVlSaOBLXlt0
jdXIZt9EtciIokHv71qAnKe4K4lkRXeSYCJ8rXrujc5tmz3oriKebpuu3Y/7bryKNY6Z6hCqma27
QFcptKFD9hDcdXMpQgJ7cA+VNRlmQbuWGWFdx8uV9Drmn9L6VGkm72KmTvQUd3LsNaskCacfhApy
nhI40eP3xA81P9bAZPfQWbaLjGcBKxJnS63GD1hJhetAAhJ/HBagObU/w/hHrjCklpVykSnPhg6c
GxsXHk5myZQjKbj7Sox2L13KY4ubDQ4PrWcMTVVy3pV/KJpuBI8tntbJDKe67d36+XU4ERszbhVn
j2E+MHtEF9yIi6b++dbs0b8yBL7p4uQTQx2JFgwLAk1MfVqQogA81jfobDxN7LivIZLReogDdpyK
4/uoOvDEybdQ5yVNrkMwzszjBulAGB48nID0LMaIZR7Hn97JhcGfjZ65cj4vCtLnHpde5vlyvzeC
fMNex2n+3WDvvscgqG5xsH99BKISPgcI8xf06b5evrNwNGXDwk8oA6WrvwNOuSh5eO6IjEgF/eeu
DmYi7P4GgT2xalG3mvn2q/+VaVlXVvOQtIuRHI5pF+zPvMVUg9GKE+l52lBdo6ShP441V6vEKOHK
vt6hu2dD4d9dnmv/XHW/2O8ZpOA8uY2cjAIrz2IFnUsRTe2sk9605cGzn0AP1SIGBA2XdQS0Lt32
GXVg+XVvVLW8gTFwdtLwW7BquGqiVdRt4fE8IqcgbYSo5QA0NXgMPyF385GXQKWVGNWg2pFXE9cA
EGUtBTtfXpF6agHIwsXbhAbL/dhgWj48+9hr++LLkEDGlQemWdntVHktXpcTOl9jM38+qFO5QKf8
0woH+FeM+waqmyaSP24lL7ra7UWqlqrma6dm/S3Var7WaPpUCQBFg1kpOUG78eOMztzbSaLDkQ68
c4ALwWtz7w1sH8sHKtbJK6tj7Jcm1Q67IaVMZGKPanwCNmdVbMDEG4WNyhChxapaY17mBwZq9tqY
/nLC6lTzdVC64jES2dcEbGEz97OZ5k+HaNDjQNAwgCUkw+Ml6JMKIdELgi+F1lNa2/0raHcFjsdv
2IpsoakFQYQ6f3jH1F2/Ha2jx1hwJXL5WgHI1OgP0JoZpSd3WEg+otnUfJmYw3jzjXpnxUBkDTXh
NN0payz31EfREXEOV3bJYGV6IDwGvwnEnt9Kry48aEv2jFFz+Nk0JIUzzDHp41F3kqyhB33Cw+dd
Kd7DnAI7VplRB0S3R/JbULd86s7Fv4zx5OI83r7Z7tJvB71wQHlBi+OOnafxP4NMp5eQBpOV1Yxa
eDaOYpz7SV8hqgkHBQmhimENzyjxC3o+pn7J09vNqzKgAs60qG9aZ/eYbzJWhm7gkHq4+ZGaJVuw
QtORMEuaV3vtiypuWWHneqX2bQjVuv/BUL2T3E6GFh13GB5r+yLxCRN0y9gatgXUXKJiApbe1Dol
yC70iHyKQN740zl4DPG25p7iExr/kjU0JF7w5JaHmYqbvSklnqnbsnF9gSzqsMlbaESG9MrPxmEB
mdqjU/4Azvf/lOk0K9FxSoB5HlIx2hT8bCRjzIZK+hrRfJVBMLKSdi/FKEXPx4+lns4tTQCnPDoV
b9zlciDoLGJfadRzIexb9T/qeTRPdQQVM8xyjDMixxcVZzKNKAAmbSRtE0db0RR/cr+JTT8sOcAG
Lj59YwFe1aFZhqoBSaun+5XvxnUUnctDFhkVQJgh9pscQPhPRObhGjp7lbblZ9/ScJoG7aK1YN7M
jihJeQtdi20nOjGOxN1ZPw2z4TmQvm+WlIzpLNTebIgL+xmQDtkZGbpiHXT1gLlFQVgjteK03P6F
V0FYQJZkXH0LLYdLUfJyZeRwZFtZ8/IKE1P0ut55zX1zp9xnwOsniTgaZEpM+SYz+OnKJqtJAvXx
HaAF+QIIF6RS+bhqZG9xPt5pNgr4TuJ1VaZkDCvXz4ydfV3YZGSSeniYB/6LXHppK8gueKq7F073
EU2ic61tfcQNP3/hsdEBMZQCjTH+zC/pIQL+Xh2qROAhKZC7TggmpWeM5oTewtef/mdN6QAtMfdi
bDdr59fOJoF45Awp9slA+ivWKnhRWGxph7V6uI5FiNEMRUHBa+244TBgCpszyvzGD+GZN/dJA8Yo
dqNN4APoNFPsm1fryNYw21xcOGy5fqOPOTHyBE8bTHP3JwZfRSqz9v5kg1Dn/Dqo7ykGidcJF5T4
v8GqaxP1tVwmmoXxlVFo28N698V7JJF34xMJAfiUsMggEOO03nxcwhx4PUBNkcb/aSQTcZFuaqp1
rNF/NCydHRpF7Lk8WDNbUFhdiMBHDkzMC/9eAvYYnEU+wv6u76zsCHyMyuBLVo49oZDegMb7+Mkf
JndoDBSDdk2UuHcBo0saDaT2k4ea3b6f07VoT+uRSSrP32lwXVf4Y+3UzeL2nw00vbCEM6sOYh3f
eJPDMb2Lu9m7ILT5GX5UjzMi+hb7hkwMxptyywV+WxEKEdvXr8gnZA63KT0UAzqk59qLVkMKhlQj
1XJ9QSdwzazHiJQ8C5CD07cAvO/YNK8eEOOcwJrG48md8mAlAfbySQkeCKNyL81n2nSCbBrqXTrZ
TcKdbPPAvjUoqsgfxvazNVCuizphsGjJezHNKz7GUR2zlpaTHfz6an3kGqq+6jLHZxxI1yO2SAPp
tCbHFsoSdIJGTroM8d0vpLaoEwCUk26wF592cGZajLg2DvxJt4ZhC4e014UDpFklcjzRgCAl3LM1
KjLriX/Ri3HyJZ8sR0keiT3tte2BRUu1u/eE0TtJ/Enau9gzkwjIjOeCQd094JolpSdMDa14fYoB
247VrRjPddOwlmJyFhL9WgDF3clt6m6iLrgQtsLac6y3bLNCd82K0I1gppKIQDobmqxjuyLOiQmN
qPyZvHDK50zq2ic+HZWes8UjvQyOLtoPkkW+GYDeu4JD5nGpMpmuIWmSGHEEvkqfVN2qT89bnQ8N
COCfcf8BH8Ched88i3wD1vFwQYOa+Yjl9SX8o3BJeWtuSu+zT+9PL3oUYqx4c6WyQMmvYBQ6UREs
6PdMY5JroQJowc9Mt8j7IgAr3w6d8jECNq/1neyJmw1/M0FEFxHvOhyBBHbdQ3Phcv5+grq1BnF4
uXELzYcJY5623X937rPNUQLEj4+/vCgxDQWP8gJ1vf0k+Z8aH9xR2ZbCv/S2bW5xOmpp/hok8dqv
QLU+InPNeunokNtlltjNMhr5nUAVOVUW97jwPbVkEvH5fRBxzOZ0l/j+OHGEpa/mUSFn4f5cvXVu
fpCvvXOaqQPxY1euq/Xk8fsDgajCKuusl34QV+H4gGFAT0FErFAk+lRXsB2OTCLRbyNUPdSfZJ9D
j1k1viSQ2PhhDGHH9WR4w5ZWqSXPaxgOrVKaObD9ZpwmtadZVw10u0FgSKlGTYj/jncPXm3wMtdM
ClLt9M4UlOeg+6KPYSqSI5rzwCAFSQ8XQSWmS95CsoXghJX3lVIQFzSBuC7NfjV9LMfAiOPtFqyf
9YcUtxS58v1AUEoaYHgJO1CxFK3tflzA7XX2LKXmF98NPeeDHk5PlLDFpU+9xudKUfDLKsP7PIJ1
6XSRj+EX5BPSQtl74+LW25Wrp3/v1mQoCibn88eCS2NERsqkGnVUGPiusGAwxx76xNDj42gIBIE3
99pebhNxUQ78z3MbZZ/4+5b9ca+V3xy+hR+sLr8YQ07jL4VKntIituRjkA9X2FHel6WD/iB7k/7O
p3Zc6r/g7Vg/GrK3rJLzcZg35UgcVfn5NdSWu5ElY9YvvKexC+qxtWaBSh/i0IyQUkQHxIFvk5Qv
jKgG8jgiN6FqjDkGqetCOJjjcLYZa8qMsWKyNdAyIp8uPI/nTY+y/B7ueYqoEVdKK/IHAo4jaO0p
Zd2CkG2EdSPgU808iZOrUsnUZz/PS7t9wN+zjQyVVrY+/oAwcEun+HIkqg8e/waxit/tbPEFT5dz
npk98AVWD00w1r84fZ+O8vG3qRGjPx1xof/P+2GAZAxPtRllATn5aFoXpcltgZsOHZeS9FT/hqO7
D7OnOkstc+3K9nVnmdoO/szGHjZ5PrKG9tiieGFat/NSMxJ3qvP/zv60uqN2g9HCAto2FvxkUzTT
6QxtfE0fQ2ptJa7fyUo+Pi/S+F8FnQQxzJqKXD5BuFy+r8WHFV90COL42YlfZbUnIl00iOsVjY3y
SSMIDWM4xoWFJbdrYFbP529buHbk5WH4ryuFYnRXBRd9DCT9Op/E7vIbxQbSc2RY7pkvqKnIJfqQ
nBJuiEz3jB/c7jzNOp/gPJCpHU/Z1JXZVH8v9sAmHLScDMtUF6OUGRXzQQnGtzZNdAfrFetQr1CJ
e0TMfE2DkJsWXXCqqTOKPs7RK+djZeGoIy7mmJNPXKyodvIZ9zB9rMXuLGotWVDUczbYD4biQQQU
TGk/AZGt5ZGN32wvd7OuKUED33J0zq7nZjZDzPJjsJjDJIv3TuohQIoGbo4l9GNgqTaRRbJCHh6a
LDX8OeDp/fbipQDhsddjNod671HuAaq6rAg1Qs6XJ890COxR1W+w+KLYn+yFd0z45VAXgQHIsQBS
3qtyRISpgp+4R8GJndfA0LPllFbVjZoxEKayp9CgbGIJNUtAEhKU23C6dm1Fmmb1Kz7P624gBJEe
2xB+dEWz5eGN1vG40AaXBVdSKCBM6yqiXH5+J8akAieNXVamzD//f03uFJ9I0IFVxz2kmA5cVNfn
cwIxYtfjKisyLj2aEy8FGadV9sEpSMoPEJBP71ocNIM7GBM/vHAAUArDqf0FMJevGJsglwqmSley
cOEUAuQXjGgDM0S55wy6bgfbk2juJJaS7BIyF/M8w+plbS7BoNl7YkWthPFdnu2xnbG8+Y6XUy8a
QH7qKYCmCxqanLqORbFAMQ3PgIuCJxSvF88Qc7t4WEr6r4fFv85Fs5HCgWsaZ2Z3MY+IsSXamw8z
mjOZbugQEjniyK7df1WvK7bo6pxZvcD9OqQWSgXAQNkjKQ5Eg0o/QC5uQluCF+fqIpWE3SbjEvFn
zxC7ZJ+2o6YocIdtC0X6nT9A67T6Glw7imYZqmlWjXnMjEBjG9TlYWM+b2EIWJuadtwYt8Ao+ILG
qpEBpFGmLIRWisslHYS2qzkAc24Y1lhAozzyYBKVRHFEgrFA2PMoD+Ar83lLiRNMwkC7vKK1ouKY
b4Uqp4A5HRJjf0HsybuEW+kxXLV0OPqtbVMG0mpMXFqxkTwIi0aHXtFTopns2U/zIRToYUdl53bp
0uX+I/BRidTxKosjZ5xcs4kMQq7bWjdd+UMoYVbAtZu0mnATSeu0YGctRvEE9aw/eJuauTJj5vDd
zQV87I+dRJoDx6pjIYD6jQiD3yVH6q6HkY6r/Q513x4ISxvWs96dOkt+DBH3r2isHCrmNYO2zeuw
ahmLKK9azVdllTdlhf7yGSZ0GdmqS3i+bqHkdTRglcLisoz8SE6Na/PXZEixVz7kDhYrUnp8zJ1x
BYDXoafry8HkO0Y9yxPJWWCT4DinLjPTwzZZwt3dXErIpzQMyE2G9C/LPDU0pJSGWJ2REXXvi+3o
emyXKrUf6rJbdaYHXNYrvTZBEXYjUkUBbdQpiYSnzxHTIqKRCQz3UUzVhJMLs4sqjgDoy6duzaKJ
9MwUH+d2Ymb2540PNpEoz/Xa2eBBxXdpO+NDFhybqLmWJvV/E6hkBnOuElL8WlqX9T3nj3S88mud
+Kbn0QmDHJseKBBX8ohn+Jr+EgoKl2DiT/ZryXHEIBRNpjno1T8bCrbj+ESLvmydhH4ALXrR3Vv0
OgT84I3nzL+m161NjUyFf00fTROJK8DELzu4WuTTvKgcDNxtZ9H62SSfB+9MlZpIzPHeFMHvULW+
BI8/78KLZEWp4oU7iRe93CzmVTvrqPvZihz0Kn/xKZFG+VV6bsjDiSlwrP7Ae/vTvL/pfrzxcC9+
iOco914Dcb1BKMaMVw3DAWTDPeXDjjsNTW6EwJ6ZWLYNleyCtyZf9uFxu7aU3T/I2aPvV9XdbKJm
KPxy0uir4uB3LElvMY/owk72KafPa25y/N4s4zvUQyAcV3ePDM68i3pStGNgU+cfd/q5n9cIiFG8
cXvw0z8YaJkTkIGkzxLcp21maprpVYLZc+ZRUIKlfCK1FWAEtYf80Ega9YVn5xbLaIRsMtrP+t3b
7bzVJ8/xVB5WHhKPNtixKdveXDw9ovNwVEzDSbP4f76ohPpqfDsKUpkFvxN0gqriFBxwNP1ZQqeU
ZV1VxHvJ9Ed/GSwzNEvCZnYuQ6XVjPXPsn7k8J1C1E+voa3hy8fygNFKbWFlXlQsOdZJCErbJ/gk
1yxMJWO0JziIu3vWK8A5URH2LCmFcQ1VOEZ+irSE5F6FGIQwd9kI5xCBwAJpKhjl6ij9HfepH2Gl
Ucmkcg/pidaU9h8QM3DJb+37DDd+dBiVM3A//5Df/iKUDup7Pic8v/ng4KK+9uSXhrlE1Umeo9Tt
ykjK3Hoasr74VEAyLZgcvQYRbe+5dbIVNUY8nZa6H4x8JcbG+CbbTLnz0FbLNbRcRN8IexqER3aM
aJlNsCMeUzj2NVxArzSOuo+GVmxV7bbkNSKwSdSf+lFyrQJBsvSvhhsMJxeQRnReOaqk8YEQMIwP
J1UBq4GewhXmBXqWnIFmuGuPEBpsgJ+0rgR0ICzeJmy0B3YCwMtJGAAPJDbqGPrXLJM11stuf1n2
K+4eMrvoAfeSemSoGHGYLXY9uF2FR8sa0udusNUSR4i8xGg+KJhSb+TS1PirpbhKt/AWMVzNCrHm
CzGH0pSHUHbx4lGNhazTgqonfwtOC+aDB8sfXcu+LDNsVGCWgXJ9yToNk3Prur7TBbiI8thxg1QR
bD0a2vkVTiOex/MmHQutIlW0vqyIf9TSmUer6mljMtVz6ijurQ2o/fVwIqRULMqhZpYv4KnSGcUO
NsMQd8rI3m8vS/QA4HkykY7Sc5i1h0fuF3X3HlUQDqA5UKPD17RE/3xZnnepuMznNNWA/7qLlLcl
QImCy3hcIHxfkIyKIFnXLvWRcHH5kza4yKplLDXNjuFPS7doQ4IRl2/cRwAi0eGLjNkF3/kU5mDF
H+ZZK4tFuCFr7YzP9NpAEizgI1C2mjwFCfipDxQt3qN1R60WFA6gzTwKHgqmWYRH/u5Z4ArhUeCk
yHLAo1JgErUTbgDVZJetxLdgLjrFVVew9SBpLnMrU/zVdkLeyYvyFICnhOS1HtUslX5UWd9+sTFy
RF4r/Zf1wHLBPhJ2QBIdjx/mlSw1MLbiHS1m6Nu19zhrs/aiexQ69DXY6knasrZ4LE6wK5AU0YyN
g+cr3aiWElN02yAvvLlD7d8LN7Z2j+oVy2c9+LiisaQ3K2xM+FzZMgTQ+IrHowU/PgHhbQjJOc7y
r/6aa7r2BsJawPKuGJlS0lzY4nKC8cz27c3iTC/fCBSmxGfY6AlGO70IhIHyldDJ8XKva3Ki6auD
Vn+Cn58b6lq+9xoshF4nBQlRzP8RNSOO0bfnVaC4JLgQJKXC9znznPZXzb1emaDFK6UDLgDDvdDr
DbiSJdg16K+664Otzq256+vZ2EaZ4b4m8VouyhEDifU9ohLPH1NkTSePSZD0W0l2bkbe53wPbX9N
772PD3IJKokuoUAZpAMoEXq+7IUMQyec4ncsw/B7B0e9jWDrYd0m4hOEPMEw5F8NJpKx9QLSxX6Z
fYvpOrmDnF1CBOWgVJu3fQsBFvm8a9Yzt/ZyYk/vzQnVhB0RqyngjZwNUxKM4j8Vy0+Pj7s/V9Vc
mnanHu3dGKS2OFWnKISxXPAQiy1WuDtX7tx2iYx7qOe10xnz8SNE+yMKtm9FLdCeQKtxsTEQI6qb
5s23TH5c+0puk19WdGWW9tHDqoNJyt5FKl7tSmNp1uXlB1lzOU8yIBwbbzWHyaxl2q/HHYXhfsVh
XKKou2kzbramLy4bXJ3t3RIEFdScpBTjvsY/ibpLX/acGelaFW6eygCmxaemSXeYz9e1DMJPEi5e
RcoDweIGOsRdQTg/pnPJ3Xy5w6TALVmaFswbNYkhLUhhK1tIOwBgwJKX/J5hmp2XMkyLUKiguKbk
/RH9NbSFV2BKoK78US6eCnBYjDE7x5aN53p2tfwmHVzRGA1M4z3UXQwakWftCTPmJmB5YsNoMG/X
ZQBDWI/Pih9fbNLi7UGijaWTaDLSOgWwq+leCDTm1+rFWpo+IAse1zS+2HanhuvcKh04p06DYbT/
scbfdqb/5xN4mk2NTwi9z2W98FM5NQC0R300jCepPFwxDmUD/51CI+Prrv3Brs09N/QUBlDJkyAA
4lSv0xD3AD5RhSaEja5bipzyye7UQpGJFScuy2FJdZVVpHgZDoHnzxE+q67NdD20y6euy9Tjcjrm
4fy1ouoRnJgMDKN+WR0e9qFQcDEFlxgao+ASKizG4NPhd1atcPuW9O1uKrBN5mubJrqe2haKZZ3+
ZQwvqXtya6Hihu9dKiwy5lqqWe5bCV2m9mGA/xNB/JkYfTUL0Cw4T2CQw9iiQvCz1Z70b4dgfiGO
7RQq/hflv+ozA2asdeoTr5SSax5GxxUT88BSI8d/zWkhDytyV7YuPUVz1YDsuOXtZ+2l2F4NDSfL
1rF52u/tGM+4pgf1ZggNA6+3FSLnRSdSmJEFGjMFasMnu0MMg0IvOVRW1gXIRgQC045hl9j97lzB
Q++yQRQvr9Ho8pEOho1whm8+20KIqlkPPn9ZGl/wBobSZX85B9hEcOd6t4SPlTVMljVqaojnOoba
qHR4R+NN0fu54eQGa1BPLZdI6OMFjAlIqevQiNYH91g5fVreoMyPi8EjlLuxLwCLIVlISi0QQ0kr
Otlheww7juAZ4Kbr4E0HGW44j14sgZxfC9NQJOJkf4HAyNvQpF1sIKUcNAooCFJhr1WSiqxh6SBr
kBiOBj+Fypag3Q9D57GUxrNspfe8e9ZVMzav0ktppoooqx7aiF4o05C5wKollIQgu9wL1lFmEn4D
DUOjkCbMZ+HWDqZcolJoTdZg/1JcSB+8T4TpdTJ92whvSpCydZH0B/jtZnLybkM0VOVsmm3JzEtx
4YSnJ5ML1sSvr65nOCZOGkmoXzSjhsIqGlSvPw79V2MimfEKkHVMHU8elVPbXcBHcrLCR1kTC8BW
tjZERnGfolmg8JwqaD2n9x3IQv3Hc96JqY1GBk/QcphhIrAzXoSeYJ/4YUOeeW9MWie2MlE6WQkr
DlPXf4DEzK8shq0noiSGX/EM/tnC5Ey+A2FRdby/2X+Lh2gY+rtDAjedWGEproXFiHaJ7vRmzx/3
CUXFgM4QoCHWGOlKJtRyYeNhvOeVtXcPN/+AHxvv4JHhp0pBcW8Gr7jZ791kdQ+vq3PzvnutkYNA
/mkLaUKnGfqXTA5F3eQEjko4OoKAPaQjEJyhZWKJLbN7tS5GZv5LOCiJM8MDbEy6JcVL7hxXEi8W
CtsIapEvHhUdyyTB0GLEN0gghE+VofoxYpG8Xhp6bTPatQvyK+vQwGDszDrYvD5rNmqEgVTQVozl
uhNaQItEmKRP3HhEvftCcCXQ50VPNms6HWfIFxP5Yt3p5sW/ofzhgwdbZZ3CUIJnACNMeGh00uf9
vqCrafMuT50wDU5MM4CNGC3K44HCNTGjc+VVULtyVWvVgEqYgKe/Q4/mYcDK6QV6+Ow3Ygz1e3yW
XpCA74raTHgODjiS0DV27Gkw3xHTThgojCCD2rxUWKa10lQrs6TnuGl65kGpiCh5UE5FUF5FjadA
1+BaV2WDA1gSt7jfzFS77T8qqX8ctr7wUHNnQktSNbeq/8fk24y8uaHhtOB/5JdGLFCyMkms4mB0
1r2a1P84Ov9HiFYWgQql1xDHgSh+QkbUU0xwbM2+MwJD5d2tVgsECkiD0Z0J0mOQrvM6mT+HWosc
xRnLf2u8nGm0m/2KVTmf14Uf7S21IBbMIMVKw7ptRwXq8LG6pHAp4o0z1tuOGBQjYIL3zk8o9JZO
Siw364QDBep0W4jtJ0Lk86fu2Z2osaBoXH8+6P8owRMjzsob5ZzGH9pPu76TjXYKaxUOJkgITTrD
CeO0TO2g7vyXG+SHWP1v14oiEcVxgfKhBUCIKAdfPyaz9vy3/mHBRUPg4tLZa0+5PkLNfmURiQFj
llUEJsOiJ7FzfqCu+YJz7Y+6PfQKp5WNV4JJKTl6IoA48A1OppC2Mv8NNKaY6MK/HqPdD+jri8L1
SFiDNMs8AKOzazb/ZtCOuy7IFu4gGlVB1Om9tT1EATP2W1x5Pm803JzDJ3vCybIT9av9tRnTuN89
+3Rk03Cj/Zx+ipI7bBqM3dh77eZ3kP/bC8M82S8r2EcLbLsDrnQ2U4eT0Wwjs4U5Rhcpn+qDdF9n
8xgOZV8eld+0DGFF8RLQnHwJnRGnKgQOuMNCdvzD/XQ29sNxBZEnZfUbNJYFRm0PgjnZ7H7wOwsE
t+elTapsvEJLDtR9Wju6IB4LZ3Uq7Ya1Y2iDQpTAC/Bknel3LRys5aPrDBzxbfCEwCMvWubEYhl0
CilzaTSDlSmrsNastW2L0JRZEbJy2Qj2rOKSk09uPLVfzZTrgk97VI0iO/RDc9katmGDO+HcBK3g
kH4oa+VfViGAKJavj4/XDn83gW6u9KYCYfpv+301xDSgTVsUR3O+u/mGcFalq8l027ojjUQVZKnQ
y7l3/ENadharmbMCG6OGjqjX+o/niWR5G5e7u3tJ84vislBJjxiW0FxD1HUcXLMAyg/XvUaGSjHp
5PYUkgjbOmyyQwG0iZVRUII+l9uR4RkHBcSUvBePGsqrzIIE6mtMReCR1NqfG1UUEW+f71/MEp9g
V9vFjn6lXJbZO+LrKKGzua9vyh5ZOCxZ3YH2tuYGZG+oLagodiia7adVLGd7AsjTXi6s27b/SYRs
698U9RVm/QZNNZuutCDdOe+RtOBMBJteyxEziKwbG4WO9NK2tIS9pDNFgkK5SporarCU2Vlxirv0
z+Cp417/GEIco/r4aGXQGRfUutLu2EF+qur4wY8QmCcOjC0ort79YGT5cK1JRfJnCJRuGxtZaKRw
sOwgwqNyk0VAaTaNCTyDWZCT6E3ShlC1DzWCmfrGeLLrU/5xhUEkJt/1mhPc1G0TNgtW54aothXL
A7wBEddzIxaq1A+fSfUy8RlamcWcZNW06gs59mF4Fe0saT8wt4wEQIXd+MnmRwJc9gAUfvHrT68/
VIEvjuAdy1M9ZrPk/nziv3S/N83ScVaYndtlaUqYSufFyuRDrLdKAdBVhy1ZaR4D01eRPJFpVOr0
nSLt6gvkROyK8iVWMPtni1gwKBfgmkbZXuqlzbEk7K/r2sn2ELx+3zM1w9EYC/JPCB8hWC4Dmz/8
ZV+Dg7DpsNU0hx00r1926pIJ9cASXUQfh+1UJo/DyTruPGAQlbGOSZVUe28ZopKCbuu3L1RWt90a
AYR7ObTacQKnxra2T89wI5WCZ8aPdDesDafisvLrNLgo8A02sRIwgEULYjrV4mKajFBMi2hT4zMf
QLM0fS4tdcXN9G2xEL5KiDLaF7LcIWOn1zAfly1SA6mmkSP79vfap7ue8Dk10j56R7b6KF07rzJ9
ml2HXkMOoBQLLu7FqqcIuqDS5rwlSVRkXsnIacFqv0isduBLb7HAwcadrd+kumxoOw3VjO56gx3a
1tBPIxbqeJj0Nf6+xj72QM+9mfe9wurCnkV8TpILygy5a5xRCxNlp9p7zKswGBGmBCRI+VLLKuqF
MriPNLVOGwZNf17gU8kcRsqAjUcndeeojOQfJnNdqV9ncEciLwr9xDRN6Bf3HBf9QKK6M3ZsaGOx
setmlq8MFeFd61CH/+LE689Y8O/oA2oR0ipkaSbgDPr7xR448QvRwYHtc2zablhCSfE/Os+SaO4X
wL1Osg5wLhJnuFHAhmeezNW1dd+i8NA5oMw3QEj71+RLVLDdnZIqRPEFDWeUP6YGqlsvaAOub5DG
fQL1FJmbrPEp6dg7POofI/VKKbQ/sEgjFcCRVfJnVY8q7o3lZW24yMzpiwTo7OKcHVhViErrCtFT
hyBC2Vjfdp7dbATSzbXIR+D2tmntN9IQ+CS2M159imdMH8/zNeao7FD563Cfrx8+OqLNfOPJ8Wai
zzd/YvY4baTMYKbtDj88qG2iC7UiS4zz1MSaBb7kyZncQqUdphNfMdVhDFZuNnYPPb65zgajQILB
v9NImu+nyOygTRkhG3o4qaFBW4cd/ZxCNDO2RWk/CYHcnAVZyC0UQkcPNxYS+fQuNr98v/BAj0GS
LnequbvaRaYmLeIfDNKXN3+vHd0rBRgeFWXA2F/CoH6huJ1+cJvB22bmMF8tUpx/qWKlB6ADpYhU
Lug5s+4yaxhRel8GkMVt4vvQ4I4qhpLzjuvuclOBt9cK2k5hAtZX4mN3wp7eexWWHYh/7BiPMR24
YnxCBDFLSYY/nJ6PqNzht/N6vd9wdgz13y20wzugZg9jwJHNXHxFCslERSuHmZCLs8xr4SUxFusR
trOMiSt7gXVxCzMgPaY7eBfV6oY4T0/C9SJZRF3Lcu8ca8VkoCR19y6VcFP5DwD2DhyYJyUrtuar
/+B46Y/r9NOF2BOm0ydG3Pjrexkvlrf2IuFoQeqIQxEwqwyjn36vjZfMzJ/9xUl2KZQphs9pEsO1
uJlOm7ELEtRQhzBoRDG6w+5rxvXMq7GNRW23GWEn4qP0bKp9vZ7QwOgFSLI1iWvxXcg9pxZ0nwJn
7+DwjExWtfRqJViL+NpXWanywyg16HTsgwUxzehwCHkIMbYafeQjtZvrAWjSvO4cMZPFKZ0GoaB3
vhmQLoyKWdjHd9u9p0RRm3nxwCM7bp5+fss+lN5+oDeroI7c3+p/kh35TKr0XExP1T2whyEM7W5I
Cae2kb4KWSdp5elt99Z8xSccvlUdO4AKd4aO9RGtcQXQ5FWnW2HSPdP/wDevQU4gm0rzpv6gwv4G
8jqqP+eCIGZdgXsid1gMImcQeE+6Va2khSkEPicgIGi12c4TIB4Vut6SOUE17O4UU2CeHTWYu30h
F6Hlweq1NWX7RdjTJOP4PcbwKBd+lghkw7dNly6PWxM8WhQHOnHUQidSW71hyp0pYbf6mVO8zR8/
CR90USoF8nntpMmnPpdrQJ59vd4NA5VNen997OCJv6bfej00MA0fXmvkwCCFMQnIUjcGvUoNmNtU
2fnT/YbKCpa2yPe+TOPZS64HPVlBkVyoabFlZBFg+4bxlsdgdobVmsubdOYVeMBNP499iDB07Pi7
a0nz9jxlXnx/nOosud8G4ovEZMpFfBswfmjY5jSWF1uvEAeaZDlsQcieNFjbhUlRNcO3rN/tox8A
OshcHDy+6hFzxdomab3Ja+LUQBizzYL7FWGKGlimaIU8njd7aGO7CUFtEaY/FzLCEKxBCIuiJ8nm
FK41oQR7PsURk54PJ+g9jjrnX11rGar8Y2lnpyGYyjxgoLF8X7f8HebkBiu4aF4JMtPWXWrOCL/4
tadBWcXciPeKXuw+SitucjdJNsjI7uz/epdT2RyueOgMlL3IIVGGurBNBFEUsTl9tb0EvFRFDvZe
Ynr+F6J4kzdodG+yjlfzfAv98PwhXOTn9wmlX2XB3uwuxKur1mn7H7zYPViL61XbQeincWAFbspC
1CWBBWfvrimpAJccgiKR4xTD6ywfE54zibB0C7BvU0m6Hv2fcPEApV8HQ4MrgaxVo1U9uQEepe63
bUZxlB5+p8r+Con4V3QV3g/Oo0++bNEOriFTyVh8OJJkLVp7hZWJXwvYHAPA2MhiTezT2EVHX/L7
rlT8//ActA8nxysosLoUxzR5DIo1EhUp8vvAww3s1uc+M7D1dc4GdFRd4Qp8N9pWWl3EfNxEsOVQ
M8la6f6eopVaRn+zzagQe60ODDhWsYLAUIH9sC6lDU5hQGozWZS1eDlVbke4zkpKqEscv07xt8Ms
jU1YFUr8Wq/SWTdrOjABdNt3eQF7L4CiT2c9MKeeiySGxcUx1Z0hQZdTdpwPMkGe8saCgCrkVOOp
DPAjmoS6VHp8w72+X19m7McLNKJalJ4Ady6lqpduGb2kG2QVt07FwzZS+mrxgr0I4LH6xCmdihjs
L44bltLLKFWiUFfLsNh2mnyBCi42CLRY6hJlWTs4s0+IhwTSHZSKSFbAEeQq4QDJQWRdWb/22d1z
KF+mU2Fk26nsIGOUKVRsVY1y9EOdcLnYuuaL6GZ3pRxoTe3EAgEPi97OS7SfGhw5o+dLE4HMJw5J
U6JVcxMyeuz1hu45TiLvQFsnPl5Jn0waaafI6YjGwWr4nSjoiyWyBUAdOEOIlaBxDsak5fjsa8rW
BBk3XDHgIH5+BPjU7R7x6a4opA1sUOsu7DlylOGUPPepWpScRrUwmy3Y9jeqoxdE6lwHHERbszLt
jzKPUEQc6HL+K0S8kesVJT+moQf9yv53uJJeOCmTfvbDp4y2STSPF+zPOJHGbukR3x9W68ZNc0Hj
PDAtBZEveam415XQk1s3XjWa5ug4TOLF7BNE5MfrZQ9HYIBaDqKxxD7pQoo12j1s824wZI3pk7pR
ubALUFzrpSRT0jqgj3nRRw/Y8y+4k8zxXKx8l06Utq3uSAL/EpU5qmYKRWx91s+qjufW+USIz2Nm
9JujKPOXMhfEwohZ/reEHKMOKpf6YoaDZYITZXQdZ14V1fb9Ykdf9nDo4kTpiogSN16YnNfBgez4
gXdPvXYg6yJDBb2Mrg0v++h/71C8VSzKPrl+l/LeNQJv6TBJgW8UXfIyVQCISHTsg9bhBzJkJmd6
yPD/KaO2Aozg0fQxDfNa0ROy0kTkAut0hXDqoso5cgUGil53j0/KEje4V4kSGE4ovlK2th+GYTPW
tzJdZhiWmNaDFkvC5H01Q/ehYe6FnszbAJNJrYb3FU8Rok07lYkO1LX8KxnSMGHLoHbd9fVgZPGo
Bvr0vACTpFWGZ0la5UIke57uTrwt+kr7LHt7bEQ+kvBosl4lfKwuz0fj8YSBvFCEUb5hZTfvr5f5
MtgwswgnbFMUpZQWS8DnkMW3EAmw1JE+2QMxyJRlHs+f9vOvYWkUbC8/9ch2sYEBiKNNCRI1uH0m
aVraXuZkf0yBaqmc71BdsCGyuxNVLXPI+J6mbNrKE4KasFBRkE+KF3er0Net8FG1Ufm72XsusMSu
UGZ1sdTrkC8yRlTH24KPtruxFGjmnwUHAkFGAYNTReGRZj62I0jB/nwH+VZYwKJXxaF13585qeTS
D/YTKALAcZrsHcAbjm+ZjMn6ZjbhV0tmqSDBgblUpVVSYsFwC2z1x/ModwusOJrHSIurRVDL4Euw
Lsgox/0GuoXc6WzrSbB1wvbsOBXW/8VhIEYbzm0+R+YlI8h7N3v8mGuFhf/twUfonHV1bZs67upG
C/tk/11ThWBR0WqvuEfEDtS3vouVglBDQDCn1bwmdPaktxhYCaAOrw4RaC20iMjU63NW5W5b3wHu
gW0SxDcSKORDEIOEpHfiMSUbMxVZGDB8bfYrBrHKmGjRZuFAzvr6u+OII0suNihwy7WqTZHMH4gF
UbzqJSyPYC1Hkw0dqoWWLPs5hZubZDaqqQY7MQVEUm2JhdT1SNac3wr4Yt1GLRxYl8i22G0mMqy/
BAoo/sdT1OH7FPBxo4KnkkA1wNkolxZsiFyLd4Jpz9ScqvpQZvnwcvPA3rSLevmEJjLO3OqBV1ic
kaG0EzDFTEslKARVIq5D0EZDQHVLpnAByiPub2+cVpLlmlmXvfD0zQp0Z/Esdrceeq8iW/R8CA8q
b7t5EIlyaaMqA77TwNupLKLIDcl42yjSFBSB5y/SU7nTX9raSZoBvJlz1NR0HNi76Ey3laV8+FY4
cfdUsNynp3j8uesw3NjAE91qZ0arYAP2jiw7DqXaXPgdu0JKHmxivNB8kMw9s1SuIQ4NdZ/Xhz4w
DU4q6y6cWfavPlxZgaY3nHJo22yotM1JDCmoXHH4B1ozmQfysjIUTn/131+2ZK+o5uG11WSV6oZ4
pLULfdwp8yCNvCgV1rMoijnK/6rIjbJQbxBh8Mv1c2G7H6I9SFKQdpwMPiT0pWNhe1foXpdPQIZr
k6rCvWTEOEzYxwylGqCWovcgY524cwQ4cZBA7cLZ/k44TtHGiqlFE2JDU59HDa/ofC3xrDg4rRLT
MvBVYwSF1QdUFd9KIg5/xm7GLXJJxeukGzkhzkkrofBgtUKvZf+PMSfLiaoCzKoHYkbKvyEDxVTz
bcpWheRW6DavL7z/CBuIVBSQWfGIMFRXRXkiMBiwnS5DM9/kKLIAIJGO9xnA0SGK5bzFkYLmyDwB
3vFiKwqhZ5yGtu2ctxRk3axz4JbBYHXe3138eR3O+cYXihxEQLLXx1Gd0IZG9O9lW/jtp9ANA1Xb
GPECJ5CUwLYl415WFY6nZdjHPYJYy7TXBG7UzqEEpq0/+uP61C/z4jg8vRtVzv5JVPqf0QnBVvJy
Yo7vUscDa/fzSasFS8esZcSVC36DniCHPXhwfYh1TvIIXoO8VUFYHu55WKAx+1q5C3ZrzPZ9CauZ
mfQdpUuaJvdrLuKsvj8zYhNgo1ThLPfRBb59mlQ/nknCcxv6nJIJ61wDU+ux1UDMVboepJxH3FAY
YIOvkhrT67tQuMIYYNW+R9Ps3J3MehXx6ZYUCXgSr0KpxgutGst1xVIgNToxo9eptUQLJeQPG+Au
o92THFFDnc7/O+N1mIbSE/oPzeYXnkELzJ7NgjERzv+BJWRulh6UFRrF9D/VtV3YnqDSRY/LCwOZ
kqhXF7hTSb0/pbU5brrgSbjx2/ehbjVSb14hc+J03Z13GdKtJEE81nfmRfJeCt8UG2RkxKwS/it2
bVJ3pLuXEcf15MNT9u7p3ZqHVDOfu1Ojy4anYJXgvam0ItpGklOdF398NrC4p6evBZlehBm+fOpq
Iv2F9/6str9hmEWyZJm8IWlcwAno9CpIQ14aqVaE2u+99fvRD0gP68p2IVMnr7Bfag/AppurH+ej
ldJg11pGAf66Njd8YIG0XnjJjOTDC8uPKbNhw6NG+bQkuAoCWJJxAfpFXiUza0sszvB5hMyhoV6x
vUwMGtldX3af8vQPCfOkCKRQhvkb+4MyjS793gp/ZyEj2c7u1u87nYsUNnpNA7GdC8OxrQyouGFJ
lLOAttiGEfKr+rMZ/nlD0dKv7sGe4uF6U+Cl1jyb2jPlG0x8AN7ySTJ2XxXdos5hTK+z/QMepcSG
8HkV93hDGODD3P3q8gcDiXcBfBcu0y+3JUnnX5a8WlkQG8xYmrumEzRzOv2MXZnIuNY697ATy/Zi
kItW3xc09ZMTZgx2EHkWEZcUARE1uGtL6//zPt9piB+SANrjnUv8QFbUtAEhsBH9i5hjacANx8co
OWLDO+5KkR/FsygnKVSxauLnRzliOE1ED7y8ZqMuKl1P32rK52u9HwY1BJNPSmdJ+FIC3tmSKCt/
+3yp5GmGplh1bFk5i3MveRCivHWceqxG+OFAPEq0LuQhJ/ev8GmLGGsAzbGTAm1YlGY0NJ0cyUmM
sYm1RsJV0Kdii6p+Kw1W4GRRLb21/fMfBn9QB77N9yPu0Wxe2ROFoCEeLGcK2+LUCEUmsuEdh5jg
bUXkr+ytrwQOsvQxyG1y4OleLJfY6IbzDmHpRXM9vukRQ9Yx3BLU6egnnqeuMvHMDh+sFpdt3xHt
a+WPFm0rJUbwiTaqMdaTex3cjQ/dJcxC5gKQyPutQfAVxJkjd3klrzIQccaiOjpQYkDGkTTOThMS
Y3zeN5uWb1RYCZyBrEi+yGaU3KoK82cQ2GAEF9xjao9Qamjv2GUyLAUU+l4YOSH8eN0LVhE2F2Js
WNuQB/bGxAkjg9EDHQutY9GwtGR+bga6RsNtNlq7o0MMTTBZe92/CnR4aubW/JT3y73uFTxJDe+a
szTZ1zbJlebs9UtvcPkBcoIPnrsu+9KQ536o5hAn1Glh9I3FpH7rHUrMp6tVj6/fFGrZBuEMFSFy
fjl5gdmJWjAKlWMHcPWV0QOg5BTElb2WHvejxRChLhZYQSN6PBZQ+oW31fELRf/ai6cWXm9eNawU
mMN2LqOMbXhsE57YWvBRTQFMJtqK8DMc0YgPLdG87EwZJfAlwvXjLMqf+NOduK+G/m0sBEUDgNq9
v9QSNEO6g4aT7iHpCFvXGr1yiIhCS5h3u44eSIWnK67+bhINqnFb0pRMbHrt6jxPpRCBDdDw6Afu
9hugs60UowJrACRIeF0Q0Cul5a0k+LaEubL3h4VZMCb3qGhRr246dHZzhO3I7pGzTsHrbImKyMk9
3ivgGMwidF6nN72e53wdeixYEFUzpwrleGOCGTxTRjc+BhSykOvF3UQka71ItkstKO8njdOS+ofZ
OnpRaQGMmEsKeYNp5DzPfKn7UYfjJNeU4Sif00L71yzJQ9+WEDGX+aM9Gkwuvg5IsZEx7r2o2u/B
8ociypaazu3dkrmt1NRNyetheF7Pk6iWieAXlK/x5b1CgZ4jH9AS+bWrnRLfo7TMY4TP5vQ5u8uD
26YRrPzpVqaio9Wmqm63mYcaoTIHUIiXpJCJtcnmgGzlOzZyGg/nOHqqtriScF4tL+bZAej0RtZG
+p2UHEWPK0Q4eI7knXEfXZTdeNEKuQInPTuORR2X7WxJQvBd9Pg74s9KbOEd/EPknw+Vn2g4BvRv
4WfVVspj6SQGShHiBNsB4eBGGXDF54iW6mA8g80UBGEJvmIMiYkErBFhy9WYYAUyZvid6HWFJaE7
gMmFrGRxTdLq6ruF2w/yJ68MLq1kKNaa2t04Y+2/BpehHWiBH8QiO94Q+gtgZr9v4ZL1ge76L6VX
QAsMUx9dAiBo+w2O3T9INdS4LER1xfgCovqzZlFuRanqQIyobdJN8S8TFSPdjkJUTk8WIILQsOuo
EscQc/Y7xj0FECzDGQlajrpi19QC2GaIZWgTShDHWoVc0GH6cpZ1wj5j2fjKFGPoOBjlTjOshn2C
5PSLvmDplgXKhMgSgPQPgLUYX18tmwV/QR7mzj8FzTaASRRLdmBmS1e1b7Xd++0sIRBdit24rO0u
eJXtQDCWG/kxzvnkTRBZiMeEQmXE6CPMHhW7mVimwOvpc+TnoR8Cy8PaolZV4lW3Eboi5GZAzyRd
lnDdpSIdJtpYT8fSFvYJHqlcQUh7acqb1ERBhyIGcGx5lWbUqAjclVTgERd+wHVDH14CEPyOOhZU
v6xGqb2mMCxhmWFb3hTR1lIusWDQ4MUBdeaKJ9dXfvoWDvDzhzM9w2OC0QIowD40bUw2ucQ7tcGZ
P7S6of0cOUU+ncyk6UcEbSERssyBOI46s5fuUiqdy1H3MoSsOL+XEk46NM7C1CQigT/4O1v/fIJP
WXmjCqc5AMyOF9KmiloFwg4Ei76lLN+M/oN/YPTYiY78NlkwVefzJbBMwyn8tWtlZ8hRI9r0eV9t
Fh18YHhg5g41NucXPMHmI3DWWZeN5Ygg0bigRwf2E4nYYphCLJCF5b28OcyTsY3UaIcC000PZnaU
7yMj3ikkEkUzC0pv2Me4iITnGwkNgtcYJPQVtflmvE6TGMVBu8Y5B637DwfnBuhxVrGUevwXJBJj
eZGDCfCBwuSC6rJHk3Nztf/KZWrMFLV31KJohxhfLaaflc3jfodTC2eJdjMFbdA+T23ibrOza/Ku
s2f85fwZoEq2zbgeFWHQgRwqw9ROFqJ647E5zXW6N1q33utoZFrqm0zhlYbKbOuZGgk0TUVp6Lk9
gsxKk/MC0RBDsaZX3hfDFUJWMpQZnghSIRWciGKWe1C/8NesCq+pihlt9EIfYDcVS8mlvqrR7jak
BLET9c45Hg13EZhozX+jtMb2kWQl8N5IY+0FfhLvXuQgTYAFONqR1XTuxjQ6BDPP2+QzbLXOQhij
e4STBa4aH1JbkLAskPIBx0KQUk6Rt7cYb+p0x01adXIxLLOVGLrSfnb6uwzZIyVdg4ngXVBmch1M
Is8vQqDoXGKE8L3myMbBwcXg/K1TrAX8oEU2RJVbSQ5gaVBSPeV2p2KgSrYmW9Y2n+JqT7ExWArw
jwRZBIoq77mybcRZSODEsYxeQpECZRk6oe9xaPTVwMYmurjJSb0HZLKKGSO1M85x99lBj/ZR+hJB
JayABf1UFrP0BoGMmmFdUQykxGdPFKl8bBV7ZAgX5GTFaeJt0EczYtzHTQ65iPCAnscRLTQVD8sR
rRTAiiQzEIpGV0XPlUSCtzka5IJmh/OeD3zOFVXdCVlFXyJ+HHxQoY2yn4qsianAHiFCu0vAMUrE
ze1iluZrJy2ueTh3Do/RLoFzKiTWZgbKX/VyJRBExn2k1uZLbCYhIlT+Q/T9bDTAZ41zw6s10vwB
6LIj24zlHJYubFvY8lzI6zuehb0QCPmkOU8Maj0yjwi1odyteUW5qsxarabnXqqGIejr3fQjEbcI
LKmNfonQTtV+28muGI8qTr7zpyS3KWPYvCbZYIrQX/RU+eWlELiE4RLrEwJrbMPF2r7BNlqX7qBX
k+ldPouUGXY2rjbATNQQRoiCK9bQUG+l1lGdyGAjPtYtXOl2DaQVy/DSDtf6J62TLH7yCGx/Leol
ryP/VDcS6rFwtslwMd7MiY/jW4clDrI1TqS+eA4o62c1+rxzNDFwsCu05Y/yqGrNM+wMWXLQvAgb
8v0WubHuZ8gK5z3hLrHbivJnNFoOU0LFrCosex7vJz9JA3E7fbyg7kdDsshHfVtbKe2if8yzO0tr
kwsyGXlMUsKg1iy8v5uOA/dCnU23t9N4EJm4adVqbcB+oBTColEQboWi/CijxOzC5nLLyYBNlZyk
dCymD40y/LcXXKpmhTivJOKM2vd8Og/IZz2uqeCol4XULVf53dCxOqAYFBZ7Xz+6nJ/vXX0MlR8c
/PygIjC+UqOd1qHBTHBy5hh8oBOMkBzF3Qt9SUsQV0REdLL/S0jtDsHIMV4aWX/GuQa5HVzbemx1
sFHLhFfC9jmIsda+DinwAYbHrOgAyhJDeqlJ5igZkOKeQQFni/4jUyBBBUNKPOE9qM1YrPPONKV+
vYZ/zJyGzNvZt1iO+Z6LxteCkrp1YJlb8QNmFcKYh0sctvxhHdVovnoRx/fhEvGe8Q62d18wI9Gi
Yy0XE7k3qbONEoeqly30Ubb97rFukVnxwESf7ssC+9QoCNucIWaOsF+xc8RuOOTiYr55E8qFAurq
eZ5DvIgQ5BDkUkkjJiZUXU0VLCkwQYkbsbuP1YOSDtVy40kyRtTso5gFx34fzhQY5VpueUiPkr05
dUpedMq25WZl/RTT7YgYuFYu6IZ85EQHw/vOIB3i8dH0+nEseYdFJXGS8YuDgU7O1ysXSA55n8kr
ytbyaaTWSQIe3HAVc8ZktL7HhqN19mxW8hpjwxCrjHWz6Gluarsjot7e6sxoqkf5VSOrMW/4kIsa
yukS7947uj1Ikf7inbi+sLTb6bIcSjq2njeneJmE+o7U9UBsCO4/oMbX8q5tHPt0CkBrMIMz/JxG
xcvNB3FbaA4WCZs/2aflH6cfZ/LI2woUNv5z2T3C+ohZPUWVcjp80ED67wBBzA4+FMnCYuZnX699
rEp58OR/8DCjLiRHL51T2FoMfUqFEAx/8g2Y8v0NUw7gjSLTd/xA48DAPplGOL2OB1QUwfBEGYsH
S8OlPWP4YQ+To7+Tdd8D8XsvAHc734YxSB1aqMWUHaeG8IXRLRIYMHJPK9FBR1Rf7ehNGWnc7fbw
L6Srx27talF76VX4MP2eX6K7AWreIcALSidPQdcjYZOWO+/J2poOXUZ+GJ/bVWYil9DWodveJoU3
rWpAhzHa6fhy1LFa99J80jK0TOk31Uk4akmdaQWdU5PKonmKScEshcA539MtdiX1xI4mzlygBbnm
KTVCgPW2we0aEii8Ye6+PRTq//Px3keesOn680qhBRZF7qbLosWCnqWiaB6iA6W2qsb/FszEWZ/6
0ZLBzAC0I8AghU2+dVCIomsmX01JIhpeeN+PRq0EQxNprV7T4sWqtCgwrrTRJOmlXdAbw1uz1bqW
qqJd7Anbp1gO7bcPB1nqmZQJupvfdvsIjoL45z8lYd7evooP0O1NEVAIVqASxeIIuimUZDfRjFr9
q6jVVnbQnKvlwpo9o/qSfRzdLJ+Uh+9BHjTYhRXQr+KF6apszlRNNJJlrZ/FTp4l7NxKzPBbB2fS
O84f7G8suL+KNP6+T613zoHDAGXmGMqhYmU57HIhxE2vYQNsJaB1HOl2y9IKwPikIm7j/OJx8gI7
+ALmnfDoURzT+BR8Hejz7bOhtpcwpAtYWsD5/4VJ/4/TWbSOUXpQReepXIc6ms+ldnZr76SUkRzG
NCujPnr0Fk11kiM+6306tlG+ESahyK/71vrpbbSmtbcca/zBNYgLBXmIXCDTzUyHMcN4Eko827GE
YhSYQyWLpUJ54tjFs8sVYXOsyqE8c01FugOXmbyg2CbxDVDo3u1/cGHLPz5+wCw0TVCy/NVWjLNR
jjqbAA7GUCPCXiKLD1xvK1/22cI8UUITj+Ju7F9Gsg+aAmOg0sayVIGDgxQTXrnXbJtm1c5920o1
jZYNm6Ly4eb1fodcC/gez/tVxIapILONLnEJ+e+ky6HbU7zAxwvOToosRpKsWUl4NSKrLUUeISTs
PT7CS4w6CNTBvq7mLQWNrYXKXGg2vflgAsdX1X5OkP5DGYINMGlxqmlHFdjEJRweLNYpcT2rp6rt
5xd8/WUU2enLQBJxlkQQfsdBCEDwfHRtZ3qQmHyMkOGQWNIWRawBSdvvZa/K4JQ6z04NrhgW6qby
izzOtP1dlu8XIrTma2hwXGLgeZxvOCPBKcuYsm/nWqCcBpj3ySZXbG1zLj4qWhOXT+YO/5dnhWi7
FCnEILTRnVT8p2Xq2WUWnddRLMl2rmIv6c/ysTziM/PGWwfc2asCmeW9+TVYkrbrItYsJvkAHBG+
onp71cPTTW4dQ4PuqFfVbR3aAO+vmjk68nLtS7QJy+cUo12JptyFW8BNLLYzi8g3TamhccSYXVJT
CsmYv3IvxGGoyNP+ly9YLkMDGhuVFkDbuof5sXa678+5N1iKox4hUaFR+NV6aFpTZtwIhU+2RfBL
2khk66Ck15n3rfBgAekBKt13/JjCt05DDxRpm7Tk/dU0mW//DPFkOQK+Gd/fC/S4A7r0xdFsmPrs
NJFmIKF3sWhjw5ecdIrHhgkUUfhZopeZp3UahYwBq+uYnVDXkOyPM1ym2NQhGQ/CPqkKokN4Cnpc
YQtCieHj6RQtM4vTPkvjLho6B1S6JotnwFwGJO5BtKXtkwQkhxi4RQbqjzyg51DyiSbpX6/Q17Wm
vaQe68FdL1cKPPNJBXEOcuETjSRngtGW+zO6lvbQDc9RuNnk/CtteVCJgmLRCj/OgBtua1fcmqEw
5bwPkkTzY7evFK0bIPz/4ip81i2sTF8v38coRxQqSf8cwOZiibP6KRifz5QRyoWzThCCburZtAhS
MSiczZoXJkEcrsEtURSNFTHDNrCmB3Ktx4wNIoJons8QtFlvQbU2oYR6TJqja2LsW0NpyEmohRvd
QruGYTBhNQH9fKKAhBdPY4hcyqATQIq0wtcc4BsN+dkz5oMiveZXP/UipNiKWy3+ijkplu3DjEte
Je58ZFqK3nb69rnOT/9s7kzjOJkMbzeYoFj9AskAIvSFCVvv18vhVyq1Iy23huORvWEwhpVY64rp
VeOqlV3dvv/CfydbOSocZsPKIOz0qUNRpNsoCTmzpUTCP4vMfe3kOB0RPfXz6Sr1OMtjUT46bA1j
1fBd44Ih9WQAT0pgVL2uHHU6yAD9yZXfnjhEEQoMXxoK/LPwrDvPm1gPJF7EI68CtPo8TP+TET3l
0fsungUzfJXOXfyVn5YoDdIyxQ5XWBJSRH6bhB7gqpJTIj2Kndh/IRgaG8ANDh5LECxsXqIlYpgH
zL+YYr31N55yLJ7622aefvf4J5mN+yWZF0gv7N2wDPx2nnzBFL5y3la5AfUj5Mezx7RtPbZ/J/Oe
xshrgTEGMdW1tM/rRh/ftM4G3toi5BGpsNoeBmSeDofBM2ygCDUBhosoT5YZsCKo0/U98PfKVF7C
PFhyzUqm2cIiMQqG9IyHJYVcvyNaIIFogAVBkqXKMP4C+itoVPsJ84Yd5AoTvG82GvKRPsfLlcLr
KCXOjVG8LPn1tadcVCXw3HTUrfw7MpUgggjLfETAfsUV7jbfrHEC201mOFJXfkoU6f011S5J/PQf
3NaCh6Y5+mecvGrkAlg8ycG+4f5iQDUXngFwbOVlwnvHWkq0coTQU7S50m9tJmIkapgnAmW6Vcau
H2m1ISugv5xRaIio0/ZIAa0c+otyw3xXKMloYUZFralsSXGLZ6v9u/RXsmkElI0KFX4o70JHv4jc
V3XfeFCB0EHdy56jsoDtdlE6u2wnTEVYq2tojbNLjn2lY4ryr2eBRWCI1URWB88xx76mAWCoufTJ
dLRBgXPL0RnJ2k0TPu47H45ktZpw3Rrh12fSySg/yfzjuNhHvxDbHl3q85t6aJ6LiwhYffKXTT78
QGkJGfqlBLU7c0kV6dJ1k9t2O06EC/FEVbz9pRJPoWEz8s8QKvu0P4cbn3FFAyepdLO30nbEQIwk
s1SLUwwnEeVfW9xOy76rgjxiYaEhXwBq+KS9RO+JoLHi4oaDnV1Vi/bpkC6I093KGrCupM7gl1xD
6158RkOxlrUcLV0Vbwd9vFm8eUk05NUr5ytpn2gMAolMhMMMrdbt4kVw4bhy2a3LrijV+YW9yGcz
yzIeaEoJkqv+NM5fmrObTD5EP3eKMFW7k/l0Kwu5R3bOOZ91bulPgLcIB9/VaC8z23+V9H47RuKs
r+lsdi2ATkwmXrHsLdlxdlXderpRjPWzJQA7TRNQORMv9rcDL3+l+EPzKV2k/CLQ3b+aqt7ugSdI
/QXK2nZFSiPVkeErBeLTBBWYFoHKTqdZObXppA2us8YJcX7DXE2NDH8RAJDwa1VmSlMrwfohOq89
guNazqVJCMkeUOINWcb4lAzpv2g54SdKcGRJk8CsHux5SBx4/RxANw0gPK2wbp46F4E/axjlmsv+
eglNeIbJYn+Wnue77mCxTCDTlzAHz+CqhUajYHJNnRUw7GBTaD5OZ0u53TVKtPZeCQzpW0kpq7fW
omC6FcCUVy5t3n/nqZGLL5L6FnGm1DYNwUtu1bpG1mT5qKOIqSwh+P6skgs7WFfAucmz3bbP8eQb
bVz5RchdlfwEwMvdo2bqCwabuTNrGHau75cySAa+7YQ0Maoss94re46lg8Xl00BvovSdXZtz0tMH
3BjGqo5Ov3u3uXOrDKBlxs8B58OyTngrseRhZNwqjOy+mkw71WKzSXlRsMUe98XzZ6qVLq2Sv+DA
dzXzlHxGbNOH1G9z8RLHSGaJAPCOwycnjL+yIcdrW2qEIn2TyEpQCgl8vy9+dfH4aJ0DSt5yn/D2
/X1tC4oqIGnuQjZuOf/3w7XxG+TKGac6haz2c9QUalW/tL6jlGAPpYJ9jbrPd7xDwfpcBMGrm8zt
Ekbpb8zJdaqZ4z62Lfb0KIqY2HUo0raEPhgrpqTD03XGDgo9Mp0qF2dI+29T86UZQeHNXT9K+fYY
IH1TKWohZT+Vymy9GLj6n1XxTn5pFunOS4R0KOnPgmizjd4rK8xr3WQSiAfYlqtdlsv9r8APqdCm
BXlJwbH9bZ3i8RACZXFV3Qnqx3EBeLPjSM0uzR7Uxz5JDbe6zkYiyzUYQMTQB2nf2ld0vR0WE84o
2NT9n6/aJbxUqTgQOW9VldYIT5dXvv7hTF8hB/Zdyl1oUlsSgyu9hxm2Qe65utDjNz9CHEEzo0lF
7e93iSUnD7lW7Va/Q6Rq2C110uxYh9dnbTRmPU+QTF6nVrDeI1LngkM2HPn14vyEyu3MKHEYGHzH
7zKl+xjSyk5KbTzESwLGzQNsjFpL83UgZ1JjPaFd7HtDjOpXd6/9qLfR4OIPQl9q7vj0JHm/ulYt
iYDnzh0L9AAGDBGnLfBOk3pY+2CaFMQn3tRZKqWVhfxoychmeiHtZUTzA2UbXhYvBTdiUlk9p1mn
lqBkrZUXOgdEHkqhsuMdVOusOxhJyp9pUY51Gaq4Kjjlt1tsYfkmBf9CoQ6ePt1HwYBppSfoDEJN
SW1fXOYnFSwrrFxE6tA41xuHCA1lr+zMzLMNBYlHvQXbPYrXNHAiXZ1qID6WiU+lMY+GRW9fjHgS
7+gKNNsiBDGOgvUKizxQtLcok7AAzQ9wcSNwy2XLYyMMAWkD06F3792nd1Qwgk5qpYQdixMg1JzG
T9zd2zy5QhK1MCcNIMCbWLSeF1Uc5a803TQfI58c6iQx2IIBPwHg6HkemwwQnkzfdUOS735ij6Ce
fgvMbqlKSbuFRqy8TznvdsEZkY993zUURHyWVbZSaeQtw4g2LVcJAwTPMW4pn/W1z8fGf2vafT9O
v+OiTJ360ilFED0KaG8prNB2JrJjRl2avA7l0fbBfzyD3qwDOrvUdRfnYfXq9zD/umo+gsGKTsLc
Uu3ukLOXq54Gr61wwaipZt8d15dh2tnSnk+R764MkCgF7yzhM52yOy52+Jdi3b+JiFhdEcvTK5rm
EPsAENvxhO/hairKoQXsVz9PtO0/NSLxPnIQHWL5FwAlpRtCgcV8MR3HsG+23jBI/ecZPY9vZ+Se
s16Mbv/rlGNzBpcHxbt7j62Bsdyu4u4l5zWibSFC436QM0kv9oi16X9HtvQl6UDXcc7h839FdcN5
YiN+9wLSSb9jR7xQXtOniHwNjE4+V2C621oMFuVDj+iiP21dyUAwYJgbTv+MLPqy/MLmBx5uUw5r
MV+F7jesRZwZerUxyU9TtMXfUg3yOpoD/pmHcJkOwBWN9mOZruLv2p6cBYS75uULaH1/soyERdLF
ibgrIfxjM+6QFfEq2ih34axdHU+/7ci8krZ9u9qNlN2SEVzUTN3YB4rrYGjiAb+JOrOrReRJJXdz
Ej8eOwQejCHPKGe+WqYccZdYMHuzapgGmrKMccxPlKm0t5x+Hb4LGW5JOBARa/9c6UeGkNh8B2yQ
ZiyN+HXP0i6vPH/SQfBjUyS8kpbwkvb2fAVJexknYmXZ0DCyAvdk2AKvHT9LcADRXSjdyEEP4DY8
W3w9BABCt0hVK4gI7yGJNCn9g+pdBtY6dnoV8n7sxzGCr4YpzV5y3NfptDtl/Xb84zSqU9Fqb2Ca
SaNrBbTFvGWHPyfTqsJ4m3kBdPO0+KpMTa8Qbcl+WBWLmlD5XL9ry5ENN7Q26nXKPebteTpdggJn
tOqnZYEkV6+5IAFRhSmbXaOpS9YK209jqlvBjzqqD1Q0GRD86Zl+x0eTBOc7L7KV1VZI/daUzjIu
waReAVc7PfY7IJ4I06WMj8JknK+lBtZntUP195V8j1ttguXePJP/UR34ajDEFvuzQfuY6yIMqOeI
yxhvj/eBMAM3Zp7iVA9wyNp0D01B1b4mVCbwavWpqZv42jT1dwyRWxILcj+YHTq3Ob2aNX0gbH2U
TQe/BWJphugwS5pVrhCUKlT8eei3XIqkGXJNWENIjTJG7HoXRwKTsx7b34qLlI/friT8v2kaFhIk
++/T9NyZ0wjVZDpz2gtOsVWHfYW5sGKf69EHaSi23QjZKnOR6iNfyOzGGRfR0m5WLXEnsulzEL2P
F7b9nTdT5XL3EQZwApX98cytaSc1YbyhTK5+F2181dNxtJishKWODgoaHnFzOH4gqXrbzF+xp1BF
5w2w799baiGiRYXMdHVaKCE8cSAVufdhTtUz2uTfhcPd0RZ65WF5Hqf9SnNCr/blfdaFpUcxAc30
Sgrpi4yZJD7qs8zLrMeY/hIKebm717mK860TPopxr4FLM7isIvOZPSU+Ai+usHCta0h9f2kXmKz9
uAuFvqoVbcWFi6CX2eQ5dfRUcLyYlBrcgBTuDvZ1Zi3jrfYjQeKVAGMOnjXjQFb2Q39c4DwtJXr9
J3qsXn1WwZ7Z5Gt/jkVcRxRmFVJAG87KtB2LCRjV8meayzw8GXk05WAg4/VtE5XZB1ShIKStJ11R
mKUEGwI8qwJha7YMMtSAPXe/JT/jPhOWexCppPZ33cXFqia6ahjN4rloO+Vmfe25jztxXmcgVQJ1
OsuX3h0CDb087qY27YppgRl/I5BTxoEXqeCRzwfe5DuVCMZw+2vdIafb8hqtYzL/+y2fBKvNv8vQ
s3hSvzYT+Kma5fmg1hKX/HnMuw6YITgUsYDDcLab4WHr03eqjEdsPqo7TSC8LsT+VegW3vt8D0xo
DuwAQZ9Co8uYJT1NnAmXQ1Z0tikRpmoEYiNrlq99dSCdtMwoEvzJgzZbz3v+irTmLBN6g3jcZ1+l
8nPvoqX/S4x5pYuBcDCFASi6dE3nAyNdzEOCaAkDbliYgEngn7b77BDxlRUB8HWjKwGlfYp1STgH
wimlrcPHEQyfPTDPweR6nkGLGOBSj3frcuZEPLrNpm9mFWuolNl7s/pKJil21LPd2utloTyNLeX6
ejErgf+dO0c6/1spEfLwTJe8mX9qxVnq27W6kI3wi5d1NTCn8EwcxcdRHsiVxtESA49iaNmZtC/l
ibEpUJ0/Xd19m0FsDhOrehZoZZOOhpXxmjIkMyc3CS3yxrPZYsKOwIBR/cv9ilRz5x2nrtxUbWTW
pI0SQNCrwarj4sLINe3u8uuhOB/NKNohIbi7W1KMhEvqRCK/demMFNC5k2OqtWb0KC+8n/RScgU3
gQaVlMWFgVfvwuhhBpiFtQeQLJFyeHQaB1TH+aMhk8Oyg8XfAeZiW/N6SznP6Bi4NlAB4NzkKwlV
RyPudO2nrXT8Lfm4IKWGiNIr6xwFNFu2AGrhlVqd5rNaO81lXkz9dXxXm7rw0vD6Kc59Dv9RWuaf
8ZIOuj82lYriwxzBCSbjoP8E9W2BmdBL5kvAFAJ6z0QKpPNe5nf5ADBYcbxRVSjZlWbfSRsitaNE
Hv9UlLn5QVktUhDAKAwaJz5o4KlhuKYSbmLg5O/EhaWtNysfK8ojZ6qIMg/OHVLypbe7C6kGpXMm
ZoyhHh8rVL8FqIT7Aw00wzMdf5XYl68g4aY1jQvhkFvtaaWX3IVKFrGeV/aI2Gzo9ahifamEwd2C
4k2L36gc4dQ5jxdLPcyjOMkPr7G8wM10eQV341aH1HTojRjU2+eAdxtfNnzsy5uyY2y5KhzcTjjq
jThWkJHpDhc5IY0cquVWv2YZKdUqR3ys42yE4nJRMxFWm5nhNRS86xnXnIrG3RFqjdu7s06sENXN
B/f4GzV3P42dyHpzcYgwYcHf1U58U+JsKKiJ+i+a9mUZ8XLTZAd06JiVoDd4Pcd8rTqyk6Bglqnn
SJ6EtudBVyT0iYyLiYur9RmI7AwhppBNmAAnojQrYlJzRvq+d4KEsDpoiqd+ghCufvw0V0V71l/r
OUKAW1NNJfhjlM1yC4yJ3TMjwKREDAmqSpb2586Y65MkYTI/5Za7JFZxci4uuWJrYccLVx9sY10Z
O5DZCL5YTi89tb4gN44Z7pU849mnDOoixEBva0B7ok+6pxWAsWm6UR0K1Ft0qYGEOKApR4YLLKsV
MyXkaz3S5f4Rtx5nTZR81/8npfRdC35hmyK+XSTj9X1ewaLbbAzzpXvNxVWCX9wthuhzF8Wagz+e
zXgj00WacSO4RipOFIuRlixtjyohEVcv7i3b+y0GbO2FKZeUalDXn894Y0185k6L1dIs/4SNEU1J
aL/eIF9Y4KSO+v1Hog7itkEb/mntffFw1mC/vrNS94qnSXhQwXLKM5NJIfHHtfwC32yTeaX++W5H
ZPHL8M1nMRgYzTPyBImQg4DD+2LlqxYom2iUcoKwLrPgbXH33mkyKBtRhbdjkGfIvcyWm0EG0/JK
rjvD6MmpxaLm2sRKjTsg+cp6kpUQGXNuuI/HkQylZ/jwDVWxHCtgv2uZwUcnhKuLzkWML65I8D6X
jgRIFnqumgmUm9V64aFQf98Ca9EDCC/sr8xrwsW/m+0rRlRS3siP3XWIabg++G289gUPc2Y0qJ1/
QA2XbmYzm8wsIk8NieThxFgPCSBDhgRpeWaXmy/hsQdUDuEYkVkMiS/N9hMQPq6Z8+7GOds8sfYP
1o97Chu/a7h1r9wOE+yZ/CC8gOwMCADEjUFt7yfzne6nXizz85VTbiLGuqvJSaxYh9lhHYPOXC4X
LxgCdAvqr6CMai5aGSXFChqV+PXnhj42dRATk4d439/+Y9aie6DprS6V12NtPteH4NXQwK3t6gPp
6Fh6btK1FvR9OVKjDh4SN6JHM8xpL0vInc4u3RfWGLF6jw28kGgz6Dhm43r2x6nIcfvOTcHYJlxg
YjLDcLrEVJdbHZ/8yI0ZEL1N6QWF23be6Sgp5t37eCbJ3f9O2p7eoykliOTlKhz8QLbhYYH+m0u4
aAKWRbW7o3VME3d0NmI4b5ZNrhlC2Ug5HquOnUFiL+xUXWOtg+QzCilzd7N/ucT+bqyfCaR+L7WZ
Ynsi2X8KVcqS7Pbm4PqU2KLQS2IRYZddYvla4CLLOaf3q2fklKVQBkyHx/AfaOv4ZvP+DRDFGejy
Pgy53CaApLKLPJlEHvPUxcksGoAGPMgUY+Wp3GSaUWAUgIs2RHp1Csz/aJEQzpbwbadHohHklGip
9oS8eN2tUSMqLCIGskhQgyTPwE0ntOgOyZRRaFIdddThJziiV7kSK03vVBQiE6TypnRSz5wCYJjC
SoEixtwOQ2V+x9xvpjE2NVg7V8xTvGLQ672d+W5KuMIln5kyGx/FJFDdAUCDj9b+S6ixjEiSEIv+
MGazMEbWwOolFfnOG6R7mVCJjY2oSooQedeJmJW0pJuttQSazKag0ZOt0sd2k5Ege5P6Hg1dA8fP
Mt/sniQla0FXYPw3A0acayqCPPUO6GqFsTXJ+dBN8isn44ebvXHlHN0nJ/8qkOcg+OxzKuz7gIfa
cGEj4LtKGVYJk6h2fKN3kFYo6TSTTVZnId6HMoyauFfyQnMXK06mrZJ4pJfm8tNZMBStMHIL6BYo
al9bXaneaCD/Q5tf5HrA/qI4cnsynE9pvCit90DqlIBmaVQQsK2KcmRK/SX4IypIBrkZJ1fvZBPI
BQj35uUOSsM7Zm3RQp2e2bpj+El8zAMXjO+Msu2lYZjrE4U0CE07jce8SzWGsXu3TbkjNuXGFvUZ
szS/TTTfxg7vJozWl8kKZwKPRaUJUlkCKsI7yvmxFnPci7sol8QwpRgUGMHCMSHMQfIawLu+5c17
eg1WKQqmNVcf25sOvQPIKmYV10IxCiqNa+Ln037k0hTAcXPFkLM7IegLhropZ5pfpPuQw23QGUyJ
r4UgTc35Dj29F+xYct/zKnG4+/cLc/BTL+GqwwnPOZM1rRF6MZgI4qB4q06VPGL2QwywbJEqgV4U
8SE4hlgvm5dp3aGIFhfJCXBl5dQBZRQGFO510gtYOTKlvxsiZeoubvttbdih0aZRRuCStYowTm08
mpqhB4wHhfNJFOAPVAqrC4EiBudmoNeFNr5W9FvUoHI+U3YKi0PSTRvSHb1w0qTJE3oyw2oPfCvD
ml7j4Xa8lajFw5riOfHzvRvOKr2pGqGTx6nVCVo7We6xmZMXZc3VNqGTf4QPR6Hfs6DG0ub93jp/
TiFZTq10mccz0+d/5Nwq8+xY2Va3hJfYSp1SBTp/JKYH6WZfPY5/DNlxgY50bjydpKoMVZqaI6LS
mGkdRlSdEvdSCqAWadDtEOKdoQnwKMMA7bXsiox4x/o+wczijpFvjyUoW94plptmCM3QacBjrJwf
mC86+knoE7LKxHLBlmG1u9DJ1j0v/89wtvAl7q4MCHC0/bgN1nAfobAOETA0KmXhqi6zPt5/bDaY
BS/cMw1RRcv2o/yf4K0GrPG6iGQ1s0cRG3SLjd6tB7w8Zt7p24eQCv4oNzWjxkI19fRJzyiGhcpo
PmoMNm/UYeQWROsUQu3yCFf3OOHeA+lAHZx4CTI9LK6myim77zAQ2AbNH9Xni1EnA/AOZVBABqbD
0zwxD+S52G5sEVZ9t168gkTWkfHXcCMNbNU93zEBur9N1cXyDDAcT5LBK3yYw+dVcJStQwVl/dO9
ktmb/uPZrilgjnM+4Md71HjlFAoZVOKjUha+PcEaIx/PdIVTbT4PYwdaR39eZpk+nMQCWQvtYvBr
1MLZwN+iutDprDYP5RhmF4TsCdgeiwQPzlzBJEfSLmbbmM1H/CTj8P63Zs+/Ezy/84gUmJG6G1lf
PuUuso6JVR/BUyaOSX8WxsSHipy0FL8owzN50jPAJNEBM3wb+IXR3HhFFRE/TQnoj1zkGOyRKFyx
eVEUAYjmEJzmYn6IzYC7m3QDH1iuBqWYDjUyJje7xKBEfQb4OfUPwW+bdHRhTun4AEMKd0UUI+0r
/t8xVkG5fY5VDXfpk2qJ8Rdp4fJjkj9Ryu18NNvSnKnROHSebaXfITaR4H6ESz6ExOtcX3kXZjFK
Wf1PBxmRWTaybCSikPPVu/06F5T6nUCWxkdKTTMGqmYZ1esDeCFkGtSwOC7NkLn3CACx7qTfcQXG
WltA8U1eb4SXXixDI/98CPriJ4uAeiYWUww3T7LGpwx7m5XQhhFkElvvsY53pEtz6YU4yvdlAe2S
zw4/1ukAXWXjYM6La4hqw/v6KPfgFgFKyfiLt/BUGTJ/5LvHCwon/Q8yj65h0y4aSgnkDL/pKSX4
q2EjgoNEOdJwKbhXkJH9CyhIH4bCqH1RppEbZV7Kroin4CTYqgZtdgdjm5x/NE6JL1jJ9H/pO+Zw
w9yGsYWtiE3MyDZm3dHUq4BCS60QvwQhA4J860f8izxQVUCOAs0TGUZcHDZFQzWl7RPzLO+DmtsK
oW65hK7zyfE4Mx07T77MKlHj7y7NRMguerG0UXrnutvVOsiDCn4GLFfuXwhJipVJm3xrAqJAq301
76uUUZFs0hP/dAQXd+iIDCQxXC+bU7RgKK32ba2ml8ORRjk4VWeF67jRrI0gRwhDeIVPjvVZx3Mg
I5SIjEGEBHupV13AFLiXXnCnLpfwlTX3bMg3j98xrhZ8Vhg5012y7ZyX0tLZEQ581gvVAC5U0zqZ
UFXZ1yf5cjY0wr/psTpDU7mBlq0NWUX5YU0okGYUd0WdUL5x4ipbKAwINLSskpVVEDx4W892PPwv
gZB/Ic5yGH4CNnz9boHTXCBuXRosGZT5+IujieAaWMNWll3gZZgfDJzTSJMqanklUbw6HOFnK+Gm
FyRtB3kC+LkvwuOTPL2TrhZGKxCQaw/LhPjH47Py/62CbwxLzSQvK2OPWvdLxHDxGBv4aPOQuT1s
A8HAZXt25gb7yaSiNDyrmfM+rMOCZgorTizP0DAt5SlZMWsH3o2HrYrUL49y1uA5ZCCP04SzCPEd
XGENYhXtiDfSimdCLcWmpUFmERirIGxqkZ+vmkSP3l8np20RGDW1jjgYs0bJLCD+gGSqdkMzNIoC
0VfDx+rxtltZnbG7GGd5nzlX9Kjy6hbhMQZNqCsUqgx3oxwsGxdLmf1i6+bNOuYeg0OsxjLKAU0x
R+S7xCvQg4zS8mloaVao0MdCrcengMhZVbVUmIg9R/AWUm5Mj35iars2fyogKVtJoECMtxfd+0lw
qK/JsnoMF8EoCnr/x45IN5E1G9fABSNUoN2X14/wpme8EC6fK6hBZKbxALYGssThJExcSKtR0YPm
n5utbFR0sGfe8ryUnbjAhKWAmpyznA9PUhoN7qOh0pQMPAqrCjcZabMXhtZbXQY2veWprvDCEUCR
rQPC1nhk4Tx55pFoYl4eYOi6LDsFgNxGwD/vMUJKj+LOKqdDQoZXWgJUzuqMbxay90+gz1120dv6
UggpsTs0ng+GmYifZStAPvEVAUTuwZmYPH7CzyCu90q6kgwuWTkubEpUjJPjq4+OsCKCegoSgIAH
shRJEU5wvojU2HI93oSJdFaICVmH4IeEsJ8JTFOJgyCG2IuSxZq9iLSSCt1yb9dwmaydeUhDV/K8
qqFH2LElBm3Xl7HtyRMiwHl06q0XlW4PHrYA9Q5kWoZbU3uyzplWrayrWHvsQ/G0o8BHvmxl1xEs
iyBe+87ZWehb7Wt1nZr20oe2kzeT/Gi+VSRvC8wm5PVJH2v/ffP9eZa5qXaaanMoeISogR9wUntK
EWt1DuJdQW1N1lSk1eUjh+16fvt+qQBi0fRnzqTq8++ZleRM+KpKPzRE495B0tijGjl87/5oYu8N
37MpLz4v5soHj3EVbVTcKqaX2nYQewmKloAMHexQNdRtQ5nc+zuiHPMv6oO91U9Z6TDEBpidIfpN
lJmVJ3S/P/D8AAf9K1/2Rbys8BQ1OtR1+a/rY7XqYO/O/6DSYW0uqBTrAX3EyufcYoBz98dFn0sn
MjpQVRNpG70P+s5OA4thvPoZgRcPGH6gdfN+lyPCUmGsnauYfu4zzdcYkH9YjzKQ0U1L4blRV00z
m7CAzkSshLfz0BooMqOij3E1qlnIHcBXvQ/4X8n8eUgRtoKCbf9rNPfe0E/2Bd5iqHS63FZzmAe0
QEQUwJ4t3mNtIwwfbmVX0Dd8AVKF0865TY9gh23rpa0YmO3GfdI0fdOYtX/1Bs6zwBj1rf+OxAo9
s80VctJ3yQRbHXIGfYkepNXCIlllfXVfYESMGkjpy6wWEwl9/BSm0CBrCs2fNcWosowEHKM+6fYC
pg0Qsgo3DJYERUWWiwQ0vko55KsRF15Nwc1qmzQIRD+AiDb+YrN/sB+8G0t3dySyE2Lu92QC12L0
8f8+S/dHuhLwjXWE8mqzjFsCiO9ggDbO+acwfMDkxR86TvPFdHuqOaOI89NT7njNkw4SLloovqwG
xj/r6jO7+pwzhsxLuojpJKt43Qq/aqFgpFhIO6ieazPwFEWNOsPDaaN1iVAyPkUGncij1wRpZrwB
8lF/7kcYEAbN1hDqcy57mk0OiOKG0RaOuQL9zdDc9A69KBerw0u/m3S+p24KZUAZ9Lue5tmZ0Ckm
/35JBVws4zSIIYNZZ7vFwTbGYcUQBgkyrHvWghTb4TWKOiOis1TxoeIUD8Qyd1/czslDQ8oSxg12
vrymgpYCw5WBE2/7iQJBX4yvhls/DhAjj21+FV3Vj45GZKUvBhVJsvOAD0f9zgmxaEtDCl91+laT
tWIX8S4yUqRjs4ZOchSFPDqabYNOzehFK0dWp4dNs1oX7DP1GbZ7FWaoNzPIojUbUY5A7+iaGdft
EsjB/LedB5mvjKOK4nU2lPLWuCGhz4tZZuNg/UnIWh6lmAgFTPtc7IwmoRIA0XDkTK8QlJsJBT7h
whbQKQnmwfU+mXYU4bhbldpz6c49DpjuNfdiaHe3Cf+/2CG5Tj7HlooHVx5mWmNMhLgejfjGDRgE
/tvE5Q2eCYX6LAEN12ISmDCbswBUdrcUBdW5k8LqhlPZJV24b1qoEBhaPimbmbh0vSFvbz60UK85
5aqz1VGF5BM6M+wc3K3U4CCHryKJFExu/zyuyIVETR42C5YaGUcoa+sDVyPf553cuJwiBjQgcGmv
LTfFy5Pi3Iiq66BMV3DGy2SBIA5ebAOqSZh5vLeLy29m70cQp9ip2p7B3vUrxm004oD0AcoiFXTC
AS+IK7yx+OHkPGX+0WnoidRsl2AF36WHyZBPSocirGs6IdCKSDbaC1rISWbGfb4UtrOQKbXQUoHQ
BmPQj/rk1dwq3fM34Dyz68p3snCfw8IBH8GnWcnZaClqfAOyZtbYyQRTwZH7XgeV/keFRW5DoAh3
b6Fnn7R0lTSy+My43f6XB7uC9UMJ4yi3UjRyaVNLMQmI7zfKSVvCPoQTTwE8cCcxBsYu8ZK1QnyL
MyW8xGm5DGGgEOp4Mz6ZC40uLe+GpX/jf75E7j+5sOA3yPsELqWUwgwK3zTeMwwyDVsTFTdPadgx
Q3vtrnfrrC9rOXEBIojxpwXYn1h0PZ1f9cbg1mvdkBqFBIw0pJmVi45h1KVLw9ezUaG4R5KtCRZC
ypH1YbqpXLnwIwDayYZaNkovVjAb+x9OgxxkxLdIRCvZkiFfRNEn916dbc3o6kghD5HOfx966Qk9
NVxydghdNeago2k2phsWkvnC1aEWazu3WXsKwSgjQ1TvxUFHK0QLXGP+t3md8HOhlNlkZ59bD0o+
r5qChdCCIUQ0yU3p1MM4CAoAoLgnUvxc9juSybp+uLEZebNImudz4RpqJU5QLgxaZAPvr+OuqIG2
7ovlotxFIZj0NEEQy/n6j5qn5nju+QmMNQwAWxcvenuFqCQQUMUT/eONYukA4657eBV3ZeIzqvbu
iltSvDNDXkl3k2IqxA+6xUnRwtB1PmkWd+8/TbB/n0DzPFyqXW0wdC7XHMYhedHG2XaLN328bxfC
64118o87hLQXLEkgL05mH/fjn/qlEKN9rPIxPlBEqAkr0Jj15XDt8EUSzcpAE8VCPov9+YTdFwud
s6pD/UXxHFDULigpUY0Ouhf54wOJhxqi5tKsF0lvgPh4DecnVdpL6CzO+9adilES3L0pfA+7GzYP
zDTSGTLGFigSZcGJKU0EHiiFyi+qB+6tKavnHkzl3hySH8l8yd4Uig7fOJv1eqtJ+9H2UT857qGc
DgJi2zEU7qttm0bGfYmM5oj/PI5JVFHVNULy4I3AUiafw6T6BSjA5fCW8EGaCoLzDoKqwtEo3Rwd
h3FdUsfQvEvbp9EgAcMLFCGRwYRd5m81dyS/RJBUg1Ue8i6P6ecLiBnld0ISAX1ikvFQs85EDMB3
mQVsTrv7ttMb8AHVnNs0u2u3lPwZrIi+x8EXYnrErzWWW+NzP4wsHtXIvFxNiVufJBYciN75QWqR
V1zcUV/CmepBZk6O9kJTVO1wciMUtICPYP0I1GiCa3vZGIqiSdvc4HQOvn+cHsVBbvfa7nTA63GY
mWrIuYviGL/+TFNWBckZSeuC19tonSEquXOUvYBAChLSm2Cru9z4U+glcfX5l3SLBRDFLvHmlXrj
XOgz/a38s0/xrGf3SIBZgMDlfgaeEETB/nh+ToKXSK3WQ/Er5WsrF626sWkmcVfiSXlsz0vZjBP8
uFdrpGthGj2yZMEYfpjdKA9WroSp3fFOAZcaYeMceu+RiMgGhkr6k25xwJslQbQ7x7cxnhWrGmjw
W+zM04acTHorNDE8Ub4wmPF2/iRLb9zuHIsBtqy5SmAYKmw6Noj9lzKFPYrIu4Fv/WRski9PdNTe
31kwYX2FH51HfDXZ6dJweWQp3as6L3IQRNZiLjr0rPmmsP6fT9UNdSPOAXpK1/uf8urLkHdJpXCb
RA0G8pcUUnI1b795LlmWct5q/USQaikaP7imaebg478WWY90l/p1R2mqa8SnHaD5DgaDTvTlI6Ex
lEHMcSSf3xJ2JoothOonq/VYu/Y0MDLl0638lpb343bfNlj8wC020uXN49+X/SIrgRwBVNKB5pmz
2gKe+e7T537KrdbVbWAX8P+7YZjWvB8+gYS06ljum7O/vtCX/vVSRoVjGa1byiGHdv5U9fGjvwiq
M7w3cQA2TQThcp+k3Gb1v6t4X6cqZGxcWSmGSFREKBXmcr4OtGqDbYn2L2mE4W8WY2i37/WU29F3
+OjDebBrXrOPH2PplhprwAOzobfq/bnyDeQNqTanwsEy5SvwuyGPeYE3dBlJaCJ4J8nFR4D07YAD
kobOX39FiqtLgb8WiedHr2bbGkkN0VuE6D6s01m16/ZkG0632+QArEvy/rjhBNA3Jr99wjs/3+mL
iw24vJ9NDlRrLPq71l8e8Vqknpu1aXT9/5fZpphMZ/WHAsc+pKPwiKPoFyxAUWqMBPtQqs+FXjnb
CDZrrpscT2gyZxbCfCSbRjMfwOK4RWx9st2s179sUBVc+kksflDkpIoX1Jr/twAH0SIoTwBbBE2S
LhNYp5Szgt1QgNK3u6rqtvpy0jZOOFsV/Z5MYUMyXk0N3bigxTlZbjXGYR8mdCHDfjH4tn1k77/W
cIgHmeSyY04X0s1ZrXgs7Xy6xijPhyTTTZ5nv/MHY2LcBOatOYoEuF5J6RxKECaQHrmXWGnaaRYt
OV/noll4hVULIhbD4GmgS4wkwbqL0Q2f1Fk2pDsWBVsVu0ZYOfoPBQpBFr6saqD4r4dV2iZlG58F
reFyEcQpBitP4ObtT8R7VjZHh6e6dSxcKocaoJuL2VRiGHMa52XzHuNc1zJVVYcf1pLakrdS0qrD
vxiaFTvshjHkGC2d0vx+IjRMLH9N8RixLnFenb0rhJhFEO5zdC1TXPyptk/IT69HrXC/K2npVf3+
rMeZAcxTg1lIgZIA/IvlPHLcO162j6+H4lwwrJDPqwFoMco5VYyYiuxDGE5L/WdXkNCDR/BfGK8Y
ZQs6EhJibMjf0z2GgsL3aMgdjyxamFnPOYG5pz+NH8GqDrNm6zSvPi6FVXajfEi/5WdbPClC/jAi
rThLDPmS1fBgUSiouyTLGkO9sUpK5wNjU5yoXHoao0Ub/5Mqlp+DG3OOmi66lzNEOBxCQat1dpyV
yS1soCY2lKqCvv45n0YRm+5aaVlSgg8Ngug3GvoGYlIwHisPiQ1nkb63tHRz2X7wWnGUGi9haa4u
jmb1rBk711W8udN7xJ2Jn7IeK8AqH2bF+vr8hJTy8EEK6B4nN7/8ODbbbNCHDTpMXIVoYksrJqsq
LPKkeappKohVAijZkr+y68LPT4vUKX13vGvpYpuHTB7FEpSItbSxCDsf/L+yVxibNGwoMhS6Uv9q
wJYooYjkPmrlLl1AAoE2WKXOYWUxetnmSBO0RinZpC9TC2JDHjqC5whPO/MQFz7AzqiKxOcQRMxt
R62qv36mwK7gcIj7QK6NRf015ZtJ8k5TR3yC+tUanyBvYmhG9LcHWGoGa5KR3NcdHBSmf3hLAFhM
W+bKk3Q3lWZBGp+uKVaWTOuo+v3rpKeaj0y/5Gn6HTa2gsEEwpr4UVlwWaYUzVe9k6Cj6d2UtMs1
zWpNKRugvNk6Ir14TI8EH+E6diZYmo29Xp1uL6J/9PTrSMi1WJQ7hq62NOVNyf/Z5pMuW3zu624C
3VJ091T+yvIBzQV0mUibBvbq1dKgvmITI0EPiGUQJ0+P2zsLPqMCL6JYrHi7Fwi6I4foyYvTx8Vv
N+4tKJ5T7zZTspNGf1VlFG4PUOG2Cy+T4fL0iBYIaThaB9t+lzeVGb/M6toFty9Kks7lcvC9Sq1e
G/gKnirwNyrEs74MSWuOPNzvxICiIOZdPqy4/qP3FbMlsD+7AwLxpd3k4GvZ0lUyayaI8FwxHlV0
SY5lP3KXqTeJ48sS+E8QJwfRBZl7RwEooNaxcTr9lyUXe5Iv5Xtl6sfG3QFJT6SeYhxW+kt9tSEu
/z0izh+vTd3H99xiUnkdeR9CYJON2pRIC/CMo/ebEuW77OgMrY2DVETG31Eb3HteVGAEhjf/B/vs
udnwvWaDHiQokOtISHs9AspSSl4+dGm9WDKeda9I6KhwrtY8TITqWd/5xDT31zMp20wmIAVSOkzz
+2SAZVFhduXRU8CF7QmCC4pglGljkuzKUmEbHuBvgwLturSBv0Ax5UyBComBC2UrTQBWc+Du0Alg
W2eXBBN9jkH/HsgaTdig91g/ynrcWIInlUFDSn/Zbgl92EHLX4UASfAzIt5VSgStjGnTcR5Bll8/
r7pCggOJOnTD1mKtVgbwQFPUt2Pp7PRsmvocf5wzupv8T+vhgqMWnTjLR/sF7lO3eAB+Y9p0Y5Ts
fBYFQAV8IETZSzOeJdl8RDZgDsZtm+4m4OScdnXcVoPvxSyNyk96XdaGjaErogKoM4squuJq7Wzb
xaV+yB1TOu7K6b/pOiybRuJG8XBil/JymfhHdO7Zv0dWp0ITN+CVhY5UdhQsSZwMDAp9fWs3+0cn
ineFEeEPoRFx+ysoQngJBjiHT++fkyfMoGXfm1+7agHGhCnB/S5I0P3T1ZW4bf28dBeAT8ypW25f
VcTS5qOXDkM1WSXmKJZ7jFS0OVAgkOuIIEx0t17CPv+DafkPwH/vl20ye/epox+2WjVCc3d1jpIR
eiGsvokiWXzOKpnBk3vqtsXMLaTq4PNjEXu+PJO4Wo/hhQrF4WxDBKkKFPLDrJoobEPlX4svKK6K
AqRIt77g6VZ3Kj9umziVtd01R1eGQ5GPotHoKvXwkcs2efydMNWt6ZbDH55JJu2DvX3QD6aEZ0jA
+QBBuVetIBqLf7dFw960cfbgRlsIGxnMi58emCV92t1dhiELp2dtRlypQltr6QIf7ZcbvuOHzzpS
FF2vDLs2RITLKP+z25klatJMYahg9+uWAUqNYCiveERY465/Ovm7/9Vfnj3HsPzpp87lev/bsD4h
HP+Qr6E9Elr8TF+1ZQK/6/SwCGxoQWaLHBT4WYnZjt1Quyzw/Ar4IBQ1ZdV0P5aIBzFZwF/NdhK7
yWgCeHK0CaLvbObtKT5RzVvoLff0hchGQ99kEB2G/kEV8QTK9lkS1zQE6OLn3Q2g2cek5VgGLTIp
vFUatXGwxU0zIxI6YTvi3z+k/hjb8vOaiVgMowF6diPrEjFlthNhTb3tcHkED6rQ/9+KTi04vX9Q
z4zYT8HSTXTsUmpSkKJmkPL6tu1sx1J5AbNDVToR3zB521ACaJSvCO7W6C/RAI2wx98KDhJwHwj+
Ii44/LbmZINJUQWVcKJ1nRCGjYnpjHaPmT7hokEXkvglM84dtzG6X3ifg735yGay9FktAFeVsQFM
B4gvafIEANkJJor3IXXy3FrRMsm5gm8JlqXpblpjeSb/CqRPPyYZrHM/xwfAFvu3o9VCo+9Q79R6
fqRuR6PnHQjpIJSD2bl2VqxeQJ+FnZoNG0olFFMdN61kCYWlBW+ldkPJBaQch9C/a35NQ/b04oLd
WsR93pZvWh4lCQakjiz9MswMaplUzX0ErCaxPhp6jjltSERF8wErDP+soP8RDRi+To1yawbECmaO
VTu+6NP6juKzCdNrvpmhn+kafZ2eqsmVtJO7vctbL8voD19pkINiXZ15Ys8zPvBTbNNjxhzRzPDi
4EbpYHMETL8VO6RtjbBEcczTR65tlmrfiS8wq2aWF2f+z9rlHeDCEc9ZywC8wDOhHHLkpeW/wmFV
RjTtlyawfCGOKQos5yARAeNlEO/KDB+g/VSmRhLSf6rWNpoHyPEJPRbmC1ZoJKaaYM8NaN/pmnSe
4KtB3K2xEqwuROPJpp9u3AHS4c2rUvytwRq1uNOe02Q9vKTD2HUdDRxOxnpkwQMIeFhOHVhYBQpF
YRUOHsvWhtOMopiDLn2B+QStAS3bF5Hq/JtZMynrb2QOnMs4w9gZ2AGvCxVgiHCaxxxbRdJROXRE
olu6O2wItaHIpXCtzGrXJlkyeNaCslTYRXg6erEBJPDYSC/RQdH2ubtbCKEupfuW1MXIB+Yu1UTv
A8j97+vO3eX8jrOH/bJBDhi+2OXGQRPm9yTXtsC3E9ojzV4qy1RSxip6kaKu+LR/zlA/8IvaCHJU
cuC3q57YwlitzYW+1S+TLnSstOWqVOE5BbTqfimXo4PLXI4qCsTDM4w3txIiM6tEaZfsAlXwZj44
UXdxKXjLSlK6oIN8aQWwAc8ASQAgvcXrHiugqAJl+3QOTbncyneOffOMqnGXTD98gMM+IEJ8BDAo
6drC6e8l61pfryTWpvqQZHBZUAQu2i3FYgQuK71ejWD4Rl9LOt2v9UBAxKFVPfoFHbn4TSXTQJps
8imVEWneqgSk4E+jeXMsqIMm6bGcswdNc5/xUJHdRKjLQj2qDHzq/X47A6qrxLZbB3PZ4dzJvBoi
M6H90cDMYudXT3P/jIfSCgRPO4I0s9LWorMkzjGDB3cbSy0mcm980DjDYTov8ndH32pjvIRKPBet
gYurtPwaa3XdggHjoBYalv3Yh6LA6WiTbro2tr3jAk51MTEs5wSd+MG0F5c/VQ6b+UiN9QQNJc5O
dR/5g281C3rYdZuh47IhMocIg/KfM6iYes9EPT5olK/Mmcb3jW89hcgONtt3EjoTi9b5YdTh20TV
pGP44dAWsnr6II+I1tYrIg8Jf/pwq1AslW/dyHDt3hk2js7OhsxZtONnhg7uxe1V4CyRTxGFAAPn
w9Svh3/4dDalOYSCNu9edqn4pc87PUEq9bZVIquabhTitoAaQvX/teXqyuXfBdgZXotWYRG0cPqU
TsFba7bOu35FT2YiKdV3Dc2P71vAnpk4wE8e5wYgZT0gX/XHwESRiIXoSGlp5tyZBA0VLnDEX5Gb
NeJf1igBKW+4N7qMRClxD5zEABXPHpdn9f5VF5uwS7u2+J4TNTWvJvMZfms3SNIppesbn6V8IKQe
0SPScSWtCoyftggMMHZSG4bLydTOcmn2QWtIxHEqlXORFIaVaVZ8xb0xidJE+UOzm/zhsc0SmgHy
ScqVthaXhhzpDzs10ysEg8dH8pGjUhctMAhlhUpzD8RfuOOd4mPBKkt+siGBJP5zhojhlC235Fd3
Z2tAGCNsqla3joBRAKY3D7SmPEXjS6XnxgTMmkl8Ly8d7bB1CAdJuHn0496MbGZsQ4iWI5ea5e6f
vKtdi3lNtgezJ3zyTJSr9wYP0ZZ5YQrTe0pypQMdPLhaJMY16F71pGLJbvj4o28oPhVfyeBvNxOX
htVtJ5UenzU3jhcjSdxdbIqH5pP77VTfeYCULmxM/0lKl29VzFKceiO6EW2AzBMeiD3tGeTj4kqo
OlKZ+bCoaSZUcqSLKvcZqZ/3OO5EZ7msBSMYKaDkmMAoP5Qd2clX8xDiTMeMC6RGM7nysGqy8hk7
LgSXS66aI8VW/eWkI5Ip2FL6pLBZNIJUp8oBXJiHLkQyA7/ZVn1MapDG8CshULrIDmiz5hG/I0xh
aTdKWFxljSUUiW38t6EvX0t/WORXqtDbzhrf6pLqRtO/guCDtYigIe32kxQowhvfQ7VC/ANptbRu
rJ2XrdCQaqB++ZQSWtKUOSCv0ShpPCxTfjd/wY++LYJtMXvycyz1sYfFGj57wv87hgOdea2Gp0zb
TAVCt6ig1buyXuEFd7bqrgUIgsPTasoZchlfBIimx1VoIUGErMsp+CT2VaPcOoASrqrEZSk6W1ku
xRKZn+Zm3GJBqL+lQqhOx7J0bXdd0hSzhRt5O4g+KBIIOO84TQnhjI53wmFx1RvOgzFzJ3wnF7Lw
EayvTYxxLiQjTq0I5S1a9abcU+uHhQS6TVIKLZf1w6GmUOHwoclgc3edlqObpBll3SuS30mCVzNH
0bcmbo/Te/b0wyCxX19+Kpv3jBLt3noBuYPipBu5e2rLXZD9R85UQT6jO6UypzHChFZbhGzMpgKt
Xnuylz4gtEkuxnmmLz1wYY0MVv2fgL/7+LViFDXOtXo62nQHo5QZsPt+GpYBwuWpE6Tj3jZPzdzs
9RoqQIOG/KqRU9tPrs94Dt3uGb8PsKHSC0nKaTxW9XMoh5p3tbWn/uUrh8fj87WD95fAc+PsRTm2
gt+jPGsMsy7Jq0JfJa+cg1I7p5XlBWy4abNsx7Rr/6sH4F1+cIoUpzQbURJdCQ9MLJEj8Ziv8unY
y/kaO8fcQ+Q9s+ZzSS8lTn4VBwunmJmNCFigQuHhM8UX9kc9qaagspoYbOZZZdg5xCQB6KXdTkRE
jsz//KxxZKib6FpCWEP3nRip1SkBbxUEHpWfEkTgEtWEStZTIDYYst2pqydOe8tIwO15Z99cqjtY
i+RHvB6scW0dh3mHSsx8H7U6NFcC9vUmKsNW4xCcGDsW7tbtQEcww8t3rxSt7JXni2tdCHLWEu7B
qMaJN9W1OwUT7VzOZ5wSYt/qHJuFQwXNfs+hI58BkBKcQ8t3tOFHMix+4nUF1+OdDXYDmv45bDwg
8Vm6MO+fKFGwCWy/gZg8npiMfvKHuzh3AmV9ZcKETkqkJnPxmm39Jsdiu8KN4EUObZVIz444QMd/
V3YuP5+mU8CuljSDWseC6O0uax341lkNF/R9o3Um7s0kuwPuor2QO0bVN5J4Yh70wAbuEAXFpjwB
12jvrx8sfu2jQVp6CvW3NVMgAK6VDqxc98f4K1rocPdO5iUo9JRwQgUnuhQuFovtz1OxrwTQjksD
v5BqopIhwWELQln4ED3HlBbW9p3aa1XgdD5p3K2t9K4Ft19rqGOK2dgAI9q/nc1a5IY22nx9T3Mz
e2VjQ9IUit0dVq7YJ8NoeLSeHLAc/7ZZg7wkhHnQA4tkxnrUVTjQ8t9M6WNvWUZY1ZkqjeQHUjZ+
KqrwIhpqvlfSML31/3QZzmu5Kbxo0T3R9RTxUF7wiVmMowc521XW0wJMt5rDkb99nI1UAacM6d5K
kQ1Tt3QVEGroNgzJoQvOF9K1tGSQvsH1qPMQk5Omzq2iDwk0qs8mxPHlZSY3wch1nKle5SOopGuc
ganzWvDyMOd/dwRtjGrX+zKBCZ267eIM2PBFyhli+ahzZtgsRVZyIH9vaW+YJiGVT1MnL530VoEO
g3SYpMPWGvmaF5qTElm8B91wCHoV3lGX6X3zUTJI02HZZ/yrgur9y91aYJmpEiW5ZsxOp3vfTPPr
PCZ+L9AHZvDR3VfzDHOvbCTwmvibMbqfgs8ln7e2HqvaklkEgFGloXXvIr7HtesQeoQcItW7ey70
n2HUI82rDYWdaFN+494hnqKle8adoDJJQJhh04eSo7QEBKhdQE7DWrzphP79+zU/Y313z7RREzLD
61Zd3RncfXK37OBx+9ABsdeXlR1Wo0z6Ep/N7gTbWrYg7cQPWhrbcqr+f3SjkpRAFsVEkPkcxY4/
y5fGjOX6zpugroRTYvpws1JCk+y+mH7Unj0H6WdPPMtUCK+/T7t+2wcjFbiSnnfAv3KOBhZk45BT
uS3LBorxZJTJvE3E4cH+bTOPzh/qDYP9i1hwLA860ob56420XCGhRmtB3hBji9zoONbK0lIGiSzS
HiUK7mxJVf/eoBtM7bqSIvhydGhapI7XR0RSt1H5f1uuSzdrVQwzs7GcyTqZGDw3jCEWQqBqYdPS
DNZ2tPHlbZFSC1BnD9s+IXi+zloPgaazapnava4M4GygprDNJET/e7vD86F7i3t6eW349QAvI0zl
6otZdf6Znki6SPuUTv3OV3SZ/Xq0omlurCmU65kHIarmZZU3CfZk9lrZfhu3PZ+sSDZNiHd3NAEg
2Z0VET4KF6v0Nh1/YtQLdNnm99Ioqoj11BYEvQuebqGdni1kaekDwP866NlpClTg3MJaJXBFG8VM
nj1FXhZHQNxK3DUpmMVR1nhr4WolrMT9q+et312mMpTJLFwFNhSDgdhpJ1BhXNaXw5jzKReKik12
9rbQfvfyvyMmiKp/qiG3lYnCaOiRKQZfPDi4m4jLNrzpukvAIPFSnTP9/RAZIpyTDyycbl5bPoe/
xFNwDu4pLzUJ1cGEUbEBne0gMRtRxYNRi2Ui2P5xgluRySk61ZKpyOlroHF1B+efbdUfA5/4+n+Z
Aj5k4/yZhJ0+/k0pxa91cbMc6I9BnSk77/FixpbzISDPwb9LDODt5daUOTgvxB8RgkmnZTKPr5MB
1m1Sif6iHS6VyK6HLCZAI3D9dkXXNSj/TWemHanXySxP4BBjYb5fMW2h89ggUbZtAT+JCSLoE3WE
fcLAIOKLsqOJH56TRpa1ZrmsXYEkRHTTTR05g0CM0rlXGUb6ioAl2cV6biWD+zcVtv/Zd4ERqOuT
xJXRYW5dCQPJWwHS6WoOlIfxp3Ze174oLhNpPsKitlVpjxPGEeNFjKpn6oR0OUWzEGPH5Ioghcfg
h3VBn4YidNHkJAgAqSCLa7L7wvK2elGI8sB7JYXdGIFIrU4Mp1HdeD+SaAbWh6jucxHEQzhIjSpv
EzPMtwklGoQktGXRlBhh9Fcop98EKgBNBXUrBLlrKiisj9TXHPE6tHdtF5kfKopZ2sPrIh16kHGX
ay8q3RLJDm1k2NUAWfvch+F7rT1D3E6410eYLkQeHmkzmA5eHrzN8BqmqCCl/9jRjrTTF9aLvlgT
pMH45wWYlm5KyWrF0HbZbX3TJpnbJGIbzW+YwADBCUt/SieLTEl/EqO1mjXrPjmq0vug3mVe2Wkd
epUMt2MILSZN2KBtDTnYZ04j4Ccv0atiNsMa5PjQ9E//5VutnbfdQMi+bpS0f2Q7sHy19nxkJrfr
F+4GDIivXBz1A8hxOFfuqXkt71L/f3JMtbx28rceC8l2053jSFTnUH8ooGJe56riNHlWWCYJ0UJ0
2D3DoZpxZMuSTYzISNbWoJtFMR5edzjoHmQ33lAYahZBuskaJP/VIZO/LroNW4NFovJ3heuXAquH
iRfdfV3v93dkRmyYH/caCcdi3F8cYWdp5LfMQyfIxp//nt+SU3k36C72kdOlJyrYJ5VKsil+LQ+J
/MIg9+C6xLQtkWrqswNMD9HMwrEe8Kj2Kv4utNY0p1o4PSByls180rfD7GppMMeI13I1yAYcC8QH
85Cze8O5sQiUlqUO+7zotjqdIiwxYaUSY2fY41amXUVaTqnzVw8S/orKGlxTARCBgdCl71z3W5Ie
n8ag9lI81kGp36H5gKToU4HnQrdMRjBAPnwN9t1lnukxdmoI+DNH/22y+kbNKPw2izQjzIxYcrYf
3avGu65cDCWfIC2hKXWtaehSDhcMtWLsV5l2XAfhic0G8gCy/Mr7RSyIDwWQcvcAL1rdOM4x7/Fa
9nUPkkGQtHUAxD21CgU5M7tAlW43+ws9enXxypw/HtYohm4csfE0nrRQ6Jz/U6/KWzAbC34nu6s2
/oaU6QmcF8Hv44k+DKzrMU7JQ01DhWqJO8/Mjq+cQUe6oJX3El6JnvwqqHegirgmcvJY42JzNIr8
GNsWsdcE09G1q2ACcew+Mb6kvHaF22hb+9vSoopIf4NWCKMhfskMH9zIhliDXRxUBubnbAn4pk98
VTdieD3hjdLI4GLRvNLdxPOxzFDONePCItPUohRTsKWNj6cuNACbzcpIWh3PrJQfuPWtjwbfiyBk
1zmIQcxwE1Wdp2cgTv5/MFLIPL8vFjdBOMZLrfLUE+iou5qv39pTYu5hwKjS1XwVx6bSJmhDldMf
9mzZlXYMKjQL6uuHlvnj71ByTs5wxCCvutPGhZEDcNRodQfBiPKpmhd8kFkKUiBVVoYygXydyKMi
z22r2giaIdA9acNBJtFZqBIaak9vxkGWb9luoBZtU6rFIK1PGTNfEBbFc0cx4l49x5IlhvrIme5D
PSpRRLwyLv9sZZv1eMALbYO5k1KO2DGV2Kba9sTyKnT2M3njl7vzHhuQn3qh3RdXOlHzEI8QKawP
4FcWru1nzA5pDNTQISdEQ8/W8Pjyip/MfyKBZl4hAWZFgG1ok4mgpyE2NDLuCD6kc482TZliNEzz
d0S8NaUiNGBHbJUOjoDYRN8/Wx++XOm5vKVnG0fjsjyCAU3O4Bv7tMsX01CPieOS4svuA5Tjbz7P
CVFybgL26dqfzT/5vaG/ChRUx99Fg7Hrx4Iy10IQkWVm3P0Mf5XBYITd1aUIneIruxUuS0Pv3xTd
3Na6bcHZRxutT4CkkDTEvqB1Wa1j7tnHrV0kZsLIzLdsZdxrC75bESX2+Jzzh6BSFWLPSsjdeq8+
aS87Mxgz1Hfm6jh9da3eTJm+Xa8DdbIA75ZB70Q8kyHRKRGxvW+nlQZdLSjK9mfncNqyDDVlvuFe
6nuThgjBe/26rrjb1t3cCEyo6I+M1gKsz7NgJW+LtrsYAa9Yt7qX4cw5riGBExRYtYIUQfWrOohx
ft2of9rqErfbTp2vtA6XAwz/lBydL0M3QLKQlXKmgDfDzUek0xztJhSWVokQ4TgHGnnpUvLxjdne
LUH02zr1OgW3fnFClnBmZG5o1B+2208jZEF3kb0wZqmQzvI+caBVOJIvdTC9pK2daGPbsR0Ukbtq
bFi9nw6II3Z1pxZDsO8+c2eSIwLGL1rxY0SDysZUjTqyALSWwYZipBtBs4vEyX0yBFoA0uZ5c/mG
qnHbtbov5AOJKqxPKASkh+Troe+ha/fhyGhFnOpNQarnYA2idhV4jbPRWIUYc426t3mKAis5PmzI
sqHDW2qN2RQE2bmYfHezMYl+zKj7yOyo65LNcssvnbn/qlLs56TZQLmF7J7qqkbyOsws8sspjBKT
QC3t9VaRAInNo65L4LisYt+ZQ63WYHmxI5SUlJDvdaAF33UJfMo2VyGmuBHJSejBkFrMSOx8/H96
CbUWoGNTgr2P5CEDK9ILQDXjbU+SJvbC3i2ELGtL61bKZ48e18mmkly9Cjfao86L/SZ2+eoZkbkL
UqSDKhIi/0yoaoe8/f/0jp7UYpbyJ1aobb29ua6+UokGSTIAXHO4B3Z3lU1ws/IZfPTpdf/WDYji
bY6x+Z39IsH1Kv90GkPqf2B/O6sO/mDP2K84OgR86LrMHwUGwmJVX5JIAgHXyR1Ia3SGhkFJfDN8
JxrpoUPOAlOUdwUOdXUnG1KI8V0/47eJ2LqtYFxXt3vc/ZUGQEwuUWBCVRe07elFdVZvM6IFqOmO
5maa0XorZN5at2RWrL8jEL92UVuUJXfT3Ykqt8ZYQs2kZgTxpiYtNyzKnCmfBLFbSCxzcbSQS5k/
NGSsnWM0uWsCLjaKN2tPpoyBV0V2xXlsYfE4B8vBagdAVAG4+jqlsnyKbISBMGDaMU9yPCVl/lFC
FU4hK+n37QhNi+BN67K5O18p6KBR167wez14gwKmrEUwa7eiVZ5ZHc0rMjbwYvH6HHgsmuy/HqLi
eP2jFBmjsx6DV79YUhM9l4esYFGV40cxDB58rxW+K/9FmT7NGixWy6fy25rerVlmnPNs3+ES483I
6Dffqzc+kxI/wsgmIXbkNObTZ0ALoszATkrq79OnFg6il45/R9qYWds7giqWODib0U7Ja/eJ5tyN
teGOkWssppSVcxLek2PXwFVItY6rtThl1l4KiWfZwHZpXkuHREoTy3D8I4iZF3L9mHS0oPLWc3gh
loHR/0MPvEKWlzLnWK2GV0RIIXF9K/bay1LSj0n9l/VRKBa9um1g3N6pmFf0bbmUgTj+a5ZdFnMK
L6VBpbzb3kDMgSuCnQmM6nmQFBd8NUanR75+77AAUhfKypM5krmuLU3Ojgc4jHLYrxzE9h8e/qxa
RxnLgKBI/0vss4fsmLsHOeZXMcZDPCEDAtiMbfuhSAYSPxsvBsulK6bAu/2Xvb7OMnqSYVCAX1ry
muzux3Ix8j7zWhUkvbSSnm8Mj1G7jIXeaDM0D7YAZzdYEmKlpjWvirLa79X6piUC1BSvnm5yn3M7
wRKU7hw+okOS+NpQoKlpgps9NqV1OxDh9PtlFFVxfMtVx1VIuaP2elaGzKwx1b64Uoca6yF/Waxh
8y04TG+uC9p0ITgFj/hKAD8bJ6TVPAz6w4X4SqjjYi7nA6q8TnAO+dirqycMe0porNzrL3tg2Vh2
frydd3uvHxIwhev7wPi0K5JqZpuDggA0EBobaqu6o0AJzszutECerr48E1RSYVF1JDIMoB/X3HxF
dskwJ9FJbDevBV0At1Ev4W0bIJn8XLUggzv1DwFSM/kBEmxy8C4ACWU+QRNGmvFJUZjSPUdLFFSw
oQiLqqX5xiv4S5+TAlV9l3G0LSLOF63MTcgO3Iu9DfvRo1j9owWz0xmFlTKBpwsCDMfmG8NFhlS/
Plcf90ujSEARViGP3h/EFnIdr1AfMEIDqFhcIwdphviunyI/C791IASPPY+NwvP6dsq/exdVKexy
2H97ZpGnjEqD9q/68fpvmrU0E4zBxY0BPM56cqMQK3qXFhSCLtGQriBV+2uiyS/Qk8ZzhFCp+/11
bEO/dL2EofsyPiiq4aYyXm78OgZeR7y1I2qzPAVr3mL1Kz+M2uQ1+3LhEDJXjcEoxdIFYUK2Lcod
6JSyp2qbwW4xj7zxMlJhtittxHBDy0iC6dGJpZ7TABmB1uv+kYsPZPzXlBik3iCUXPdOG8UwGTwa
OoVVcJgWICx1PI96cra/qT75rpynZbhOD6qCzRo0FiHFZCbW8mX0OrKhIa3ulJ/85rov0Fpnw5aZ
nkEHqrCn28u2luSFTYGrg4CjNmYQ1vKdl1YcN5kK6EG16rSOf6xY95ivaLoPeJo5nNJeEu5LTjQj
O1i0Dt2CJEgwW3OqLEjY7LRk/1PRxsz+I0UI+CoYe407+y1Ew2o2eJHSGYfloYlorpBdVgRiHNYq
qfOVQ5E98eqDfXfp6RggnfqD79uK0yJjzs4VHuvKyf1j8QctcddvRnrcXL7lHGHTZx/bVHeWSQlG
nue5qbl4JlhShnEVpn31iVuyvHLKxXEeb/Ht+8knMbjq6Dnf7Wa4NR7FDvFZiHk4VSbGcbKEPc7J
Zsxq9kqXoZt5qwiuOXRNTZJqxmGb4e2IhWDEFDWg4m/VqHcYP6Bx8ikSYiJyV7D0hCxmQljAr7DR
WGILLp0Nl8mwN/TCTAp7SJaEhCoSSkNz1oMXBB2QCS9J2GRoiEaWbxDBuonAvkjAombMHtvPL2an
GMwKPlZVUpuwosUMi8IOhDiKRuGRZG6X+/VjwmoKZkJD2kS9Mxesl80RjpBIeO8rtONjgo7na0Zf
6RAao/+Bq8bgaQRb9XiBaFVt1ERrU8CqYDBodIiEBHlBVqW4NnNeSziu3TBxLqGWNr0AKSgyQ8vY
mPZooMTSyIDrR+OaTYxXgtpLjgLkuvzlW6yQGDuNY37NakFb+cTPCJF1NkiWwEapWlV/zNTMAMHK
vGgULgIknVS5ByysQGNjai2gptwmX/9fB1Pv+h0FS4i68KtN6hgUsWPGdcyM0r2g1Xv3KFQsvC1c
b9omcvgs0HBODV3HrAUl696heuVLa1Rs6s+ZZQMxVGAJRYEuH/4eRNKYmo9EqcPrSy5MofLNTXCK
4eQtJCDy8k9wlkHJd5kfecjgfEvs8hs8In8NoNLF1ZQ6jgTbfbH7my79gW2aFZxBHqJigaPtqOlp
yO+oh39F0wBDK78WcWKi+Ldo56GDJSTXuLpF2yvOp4U2Xx13rbw1a3Y/fSl+NDTpFn1polxXUm1x
S6otn0V3veLtGCCoGDKcer6U6y84JRm13J6Ne8/Vk5p7y1vKfJZvCzjpvzCHR8U+w0OYOJs557Yx
z/S12a2K+Mw+wZAg8ZMv/CshYj7MYZrzIl5ExUmOpoCxWePLTQ3VVivMviEmVogYb8LK+uF6KVZ0
ChHltHqm0MLUEm1toa69/sf7y7MG5xrrqUa4e/u2eSfZMULC5WS2kGCwS2FiDz0olOppmrdMRsRX
CmtJAYckwi4b/w+iLxgp2extmwKhWUae2s4lgB3V+34WTO6dSVzxgm/Py463Aj65MqY+6sn683uI
xm/fVI7247HXAo5fQDZ5cgm90TIyn5//QmenbF9P4SVCd4o8VofRQ+JYlsNH9dbbtDfjw/hsOhIT
czD/GxETqjFHkywsOK0J6MHX5Sw4IGwyuq3lqKNzx0dnEkHJyIAdyoGVEYuUUlMBPCvAB0egFsoR
akKddDtWEjq5/g9E+6SrK995IlhrMlZ2VWbYYIoIBCaTblt6hOktDOwxmjulb0bUUYDjYWDcoivn
fcC6rAb2idBVbNnOFQsgGRYmYX7q2PPZWbDDJa9ft6JcIxG19oGEEfFSRFsa++kMQnbY+io2DDX2
C9yskeQea+3V6m8r6xoPD4VvKYksUBUCahc+QRWTX+oXGaEr3lmd0e1RCs9VvNcpHVFYuZ82Hq0o
jOW/mQB+nW4NLrdGYYnle9HB9EhvR14LyaYzOGG8q0vGeJvobuHFUqh7Jt72Nyj5rwZCIngp1cRY
/kJH20DLuCNpNytKX/VeYtt0Bv/xvu8LeBrBrG2wgrlGlQA+sKBX98eEZluSwYfghePMHP5g756p
u+dCacgQ0VdxSN1RUIN/8r3GOLGBMQQ2h+nwl8DwqJp4fu2WRgdV/avw9ujw2sh1NJkexZejMIcK
tdxIQZWpKEl2A/u7oFqcRlask2rVN9etxQ5CNUb2MQ1Lj3I0e0lSe67AG28N8bOf/cdrW/me6afc
5Cohx0G593hCj6uPkB1zh8bKW0ZTTTc6cRokvP6JqGT9xRN6pQ25wExJHIDTnlMzbVJ6yjGGNrVc
6IFeKZ8MSrqQrRdqPjOgT1FRajyWVZKT1OmmO1a7k9JP7aBoLFPhQDcoB1CXP9ipWF6F/Z7BlZOo
G8BwJN1K2myFFs8pg2Ou3/AZgYKJV3u1VJbonIOH+IpbfFar082pVdAKivqPvJ2LG9nXERt7w0qA
N1oEWun1LsekmnwLqmTm9yQBH5SdcWqHLexuwbeMGAitJR4eR7L+bS+QWVM64DCAx/eIgIDYCEWD
dVm5/8oNxiMr7eRfEeSkZCmBx5jvQCPc1slmuGQIyeX5/7POT6dM2kFFOFCNoyK76+qu/eK825Do
WPuVsKlwMkc7uVWI8YG5zGuyysIziGK+ppe6S9+r0jQKO+dlMx8mqY4XCohHIEWoC07F+RB1RwWF
Hfcky6Iwxr4B4tYdT2UwMcd8SziXeO3fn1KQK4krbquK+g/ltWHPi79nJN26b+gVzrcqktE7/5es
XRhSWaDm28LNPp4TMJ3EeVa3AhsLOiZRI1sj2l40Ou0l296MJMudYkXLXwAvOwL/kxQbBT6Iawd0
y3YdEfDC6xMcW2R/bjjAOasqSZgytO/FOyEcS/Ib7k9gXuGO8FnYq4Llmtqn5Z+q9m7Mre1lxCr3
fuUYzZ+tTXSSYdvj8s3Pm7VY+nrbwN0+gnHVfip6gmsJDYNFNPwmzC58RT2tR8S+w6XIpzI7SHBN
H8tJfEittKsFIzpWNgom9CmFdspLYTR7aczXxeTIaLTw8fzHaLzApoEI43pObwAfdCWecixvlSYO
RRx84dDn9Q9jOLQjU9sSHbPf7/uV9VMVYUw+X8R5PVZOfGuZcf8EourpmAtaXzg2T5iKemoISYOm
LG/BG8K7HheqyC7M8/apULMzfP1PbsWvOY5o4xuSvRDYfGwDgHO923UBIb6083qavB9308ektLkK
0LXiPuasr6VxXtN8PIL2LBLpWT8mHnj9VUIUsqCPxFShyj9PLrbGSYycFiMKqGw9sOn9sPVCECy0
N0DmjyLJq7h+4zj1irMcs0lqW8JCbVrU7HrR9XI0kU6/920ZtT13AeDVQygqrChGPvI0RMHcPaFY
z1VskQdHfkRKk0bNvU8Pa0WUAei8wzzotpcRF2byvHWSjVKeZwyjV4omVPZdPN2ea9FkQvqakZzv
+8QPg/F6KC0P895Lnpb3E/GcpGSL3AY96+cinCEb1B7L5rVdy+5GygynmGBDLI3aqRkSzxW09/Wg
GOlfYLmJD+lVuptCnYuDXpO4KBkv0exG3OrZbl4IcdJmv1wP4x6/WOZiCbANBJzT0eIlBLAVok6p
P034cgXjCNlpR+26I6NV1iXpD9WtbfPHwja5Pcw6b6byjrlx0N30RAoi4IvipBthDB+c6ouuj4DU
CerZHOqrAlmqtGjzo5lQbD3u3SUcwNQROljAfC3eEE50KOPs8OsXqaAGw944SJXbD2BXbWJslwlq
nG0dTKvLzBGMWgKJIVlPlNqtwnjzNwBrv3n+ktA0NRUkVp+43zzbrXfvvoUrp/HlNHGxJIbokk6P
kxPtTVTyC5R+PQ+dhjhc2AQIi5m3wySCqu5MouOIztKjp5N2em/v85VM1meq55rj8YFRj6eqCRbK
/vyf+1fHDj5VmkEkRnmN+Xaxj1nTFHbDYZVW25o+hhq4BA/y4bzxuCQDN+DV01JsTgx6SVk8wqBe
O6wi4+GjdBLrd+KjhfeKiOIAN3xQ6Td/1NJC0j2XpsyrjByM65N8MHEACkM3zvT4s94NGvvLBZ1R
k8QVqMVUTSaIpR+xiIrmJEMwVdg7Dx3yCBZNxv3k20Wri01AS8eRKm/oNGJkrmpIqCELnxR49Xa4
Zhng0VlqYWcSJ0ZVSZHiBNrpx3n+uVHuavHQJ5J2OpdvEjTTR1eL5sl4drwZNLljBLfqw2lZlhVt
LZkxHFa2srovf3X68LtlBQ84iDP2OnMiBzfcy5DE02EW4ZgoUgMjdANDOTSCK6yK29CbCgQZCY8/
etTduuULzNsPgl5Hh0HHaHjMOeHWW3Q+irvr7mAnYeda4q1kfz0ZmUsPm6rs1B/Kn1Cw7nAN4ur1
7TxoXmZ1czw4GUED0a+wfoRuLvq1bZqNjRPMj5TYVCdGtk33kcGCI9orLkMO/n5A/LI6GfTeqCwe
riDF1m3SuucL1mJ/uPZ7vVUYGN25ZuODiVQsjDYimZOPxbs4wItS13cg+2CBzYqbk8k/7lmM/zby
kkBx65yPG/7XRKQ0YCkj6cp4Bgtf2glIJzU28qacyKXY2+y+ehiNdYyas1YJmiSxECZEo0YvpO9w
U3KkPdGc9kbBaE8L0XXbaoAKd7ALfWOkxoW84NcZ9D0E8sB0luIdm9jxBx6PYqECZKlFrEIayVo/
4skA97QSXRFcyanwMx04j4RPFBm799jIAcOjOgCPx6/hwN06hcVLI/WXQ5hzUXEjKLCvWdl+N9xP
78UC68KvAnQiWs63bolAp+Gsm1fnSzsxFxf0mU2psrNjoOsV4yIXG4HLgo/j3WXIMLg4/Q150IQ5
9qQbR1SJgtOU5Cbyvz3c0Yjeic8Q4CkQepUW4Yo8ncEkFIMEuN6mDdrwv4TBNVXrvkccLf+iRnm9
zfhhb0dYUO0JiSWUtAWyU5RCVzoRHF37gEzy8+gmK18FkXt7W70QRvICeyND37jQAoxiIk9YuM5v
i027xM6EjlJnD4+2RYGy/U+aAViQ+oCnMEqvJnaV9QO3357ltJmKN/ZuflEPA+j+71zuCZHKbIb+
WhwHz7h87sDvd6LlVDXGoTJBZOcQTY11viOSov4o6JITCXl4UqiO+FE9d1V+h12Oz+20l9SByfGt
Z/AXZTlyNmn3Y47SuCKJ/qQ+SpggkmIROM8ohafoJ8FmzACpuQf/lH7MbqP9sHxVXWEVwfMTJ7oM
Gy0ZLmeIUTdceecYEaj5Duy9AEgH8S3YJJ/gPn5KlSjaZtC/CoNArZUTnLdcJksvIGryKBC5AYaC
GOp+JSXDwlKQI5Gz1gWxPu1PV3joW9ieG5c4VE+p0/899RRg2x3jtgqsEay/9tbMoHR5b44+et8P
oIR/Lm8ADIALmritxqOYwMME4n0lfFw+C15nMEpTBcx6K535ULxcS1KBRcvUJH1CMQ1uMsSO+3iU
r5reVAKkyo0Oio10Oolk7eyin7GQA/Xv9aqLiL7BSBTjrtWX6k9tUkYr5dXPd9aXqAEepe/oS3ak
SPLJreh7yXFQyFZxF4BF2seP2pBmYyBsOMzg13gHvQdKLS68rUEaMfN0s5AXavFTvJ+6j31jN6VH
i05ZizeglXCnf8Y5P+zxwQ93wMkqQw6W0offUC1LRPViWOkc7qoXcXxiZ4uzvhJKBwFpNbXISPo9
54XrCGSw2Sea8UwDM+ywuF0dS6H7VvZVBVViiqbvd+F0FGwKUvhLLV8XMHNXBXgOnj+Q80PZAAVr
DHIod9wKxgu5XQEX24dZgOLa6Uxotw88sNUrMfqYAt2fao8X8ZJnJC9UiXp/geOiUY9FB8choGpO
QcfT/myWsVO7si24bs7CkLsTlo6Nh2+nlzpctXlc0mwmSYAns7tdqxqTUNKdktey04Pc9QRPIHGw
Lw5eb30sBWlg4+AIPZbRolZGyFbCEAfCq4W1xBzF9lKXflfUqjWXQiMps9m9zjhb2mJ8kuB708KF
2DMphnTd+n/UMe62d3GYGDVDliXfm64mmYwpAkCAitG/rVd+RnmmQY3coTVnKOmakF2d0gjYAFj0
pgvyMdi19LfpA8C+5zBelSnRrxumeSvZDB54fVWWOwY01eUf1Ic1IdQzZHTecQwmdpr4vKNlamOA
4Mvj8pida7+YNIBJoskv6EExKfolw60xmy6k/0+frqFtkTVWD2oosszJe1YmLDN6LExl6jvLR0oV
vT7ANwe+O8mHDi7DR4GuTtjNp/fRPhH1JdduglHeH5xLwMx8LQqkBKhc4RNaeoTrAKSHatOibI5x
yldtdj2HZK4cO0u0bRGYGh8s135SNE84GaoOtqwNaxh/9hPGipcWd0/WhGqjfVuI1ykdlR1SdGL4
lPwZ8u8UHVWRI4uwXoi2yZQEn5Nc1OAd/JCt2GBGZgl35rr79bil2i0PKUXlpZzz1a3Tn2akEw9z
HCEDwxvJ3O7KHWtsQXZHxp8SvhsheSAcU7QSu2qrEVqJpWoCFe1cq7Z+qvsDPo0FHRinrulVniSa
ZZR9nv6TzQAbAlgYPwkUNePkjXXnsITpuZqgVtx/wbCcAwvN1nIyw8SPd6EArlYPvH9oPiA/n3Ck
nEDDN5gP0hlgOWbXYrxX9Sbae6iE/BTmdwtgrSrtWeaFG6GarD3DzmC+bMVO/IJnkbpPEpfVaCda
wTbNb5rcdvYqe2LpTwjTIQ4zxkg4Jwtv9jb9pCJWch9myM3+CIBM4VIz9fi1Ac9CmJXmKebwoE7T
BceZpV0MYpb3hvjwxaQ/Jl6GzG+imRbMPwpzBozBT3AGH50ZGIdPjQl3lVMwpmNa9/dQanz/B6fN
/8/lCvvGSVC8mKBW/U7SGt3EbasHObX9edQV3HprjYz8cgH4TU2G//IzdJV8heJlk3RnvXoA9WsZ
hjnqQXTTnA2HqgIltStZgEvRPGR/nGQ4oo8dc17GsbbOQpcvy4ltPGFFKP4Nc4HeQm7pvRzaqzDf
77I7vrraSCQINgzkxk6udtxMHo4geaZGEHhdjVCe16Jr9cl1/eAtf4fv5N5GNfyxZxXjd1lCB8jA
yq2xlLCa3X9kSSQeJDEWtgh6p0Mglj12y2hO4ZQGIpyTEjQlbUGZq2CN9JjPN9SrxUQ2cUdXtbTa
R8KtwyKoAoP4YAnHYeU2RLRkg1bE+SnmR5ouEQSWDMdG53MJZuTgMle788TFJgfhaOkQD6xyXozz
t9SFdz4DmqZtwm1YZ9wR1xcHobIWxWGMWZWg1P9AWtsl24xvPwtttvsC7KTUd/gl4le6v31kBXLI
w2VcoxvG7DgcJ8sPuV12d2Ye/bydvzHhz72v/QDUXz8g7oInhJ+Je5aLCkwum8Lb1zHDWta9W3re
lQ6NPAFEX3IUpetCkFFvsuYkW7TVHqfEXXgeBsa34r9yidXKGsGHjZR9UaQmIIycuCuiQJVPIUru
OQg1tggekx9XzJbWSgLG7rtLRn0uWa0jFUrtew6kpY7bNlUPwdibyIWRrE1BBYh+RTlSrbwvSmlb
0auBWsQOU3VT+Uvo5CeqHRL4fOu42nNLXPg7mDC+hVsk4Tp/+q290WLF8393cAU8X8L/d+rLLcHZ
lfZJ4lrlJiwhRTaIc9hAavpWUMMjspuyxfJxMDBMbT1CmiOLzmVPzPUtkMKYU66JWeFacAQqs7SD
X3xKfyYdtGboCSwR7uNF28zNS2bhhnzacj4jvifhHOVfRcQfg9VwV1jF1dHWMNdkD/yH14BrXZnz
hYpOEQfBNcIIrvgRf9uh63K8o/wANdH4hKTRFPajh55TEwKW3FJolmf8a5aSLXSNrct/il7jHC+C
2MdRrymCn4BFEZaYO9eC7A2nAGaS9HbBiODQiQwDPU41EIRiiY5VJoztZUCKvojhkloemgslHurG
VvY7mrDOXWg5yxFRB7VEMBBczrKQoTcdlGMsarg6jOa57efLB5TmphlyVa5dI+Ew62iUhmxg6AJx
NS4Jz1ZFfu0xxC2OR42kY3bXSqujrZyWBtF/GoYzpyfmTMukpUMxw9bJRiy/jQqWMviJCzX0QO8L
EQmcji1WZ14rKFKQvb7ZiJ0BNSiY/rYrluLoSF1bvucrqH6g1ZR4ypslOlahhKVhbis41r9DbKbD
vAbbSB/0ACNlV+wDLk5K5tEB7j/MiYLrXsBoKHRoyU82wOzM0laEsDlGnxKYpcRwh7A4dRy2aVzw
MuylzEnr35DvZjV4dNEY77mcSHnMNLxGckCT5EfYdYNf6/ZaKYBkJ8m5GtcBWFdYJiyy5ZqL8iLs
U2m+aI0fuqi/dLuUMbt3lC31qRYKKRoHt0mRMjQHWqu7EPAje/FvDYqeKADsCTHeAw0FZrZf+WcI
HC4IFWkbeDY7ew1uGOcr2UUHM6tLDOUy/PDM6rIPAbULO+jSwoHMW09fGR+boXSk/D12jnb+DzPe
+nmMUPrZWFWlDI1wdJmAj1j1zd3croQYFdB1+QBe70yaDuxg/VhT0bt1mJLAd6XeIDApalGXpLbp
FWK593MepavdpRqTAnSyy/+3N+r+Y0Nd3t8sN/4XI8erIJyNFgeLMz/VkBGUNewPoIdV95JtHfR5
38yUitZnLk4MloLPS3RzjI6MN/uGSuAvNDIjPXz9Oo7HyVIubw7FnuoiAyyjgvzvN2LyJrAo9ET5
dyn2X3EbknMgg9pHkoDMlDIe1h6ag81KHAOmx5WcuaxFsxMgyEj/o2GHEG4GhDrU2P9bdWp58aXM
KNePy/wrxt0nwOi/ZM9cQqlOGpg6GKdS9uC/qZ79ZJmA178AXdd6ES/sBnP0mE3N8SyOZWmeNQRD
xjd0rl8sqMJUYePYotQpmUz4RBh85mRydLbMasziY9zRGAl8yr/twT9Hd2Wm4e3raqCofeEYCuHi
D0RYf6SMuGjD6HEA44Z9YnaUeRhQfjdpRNnkq9qtclwPkeKRiukdxScrLfw2U8PUI8U0bmm9v81f
02EobbZvgLgbj47ssUzMpAt26IAra3cr9w57IaliaVIEKrRBzAAlZXhLsR9b5zkzUGmQj/zcsL45
jF8ZXSHqZ8HKY+9vsPdvyEkiOBspmTd5baIyt361SMkQ78bPpDJZlRoJWyHWuTAX9O8jimQep2X5
4w6TUSOO169WQAeE93b8djca/Sy9UcEIAOlsH181h/5GqVn3ggfYpq2hXHglYqPuEGquTp5nRdY/
FD9WHxjCUMoiU2vKG9ODfNqj9R0Z4p6A/hDdy8MBnghtAFtpx4+G9vnfrfy44ektweDWxu6D/0/Z
EOrEGcfozXRobbaHn31j+AHg+SGX9XMWhn9X5KiwmV5upphIYUr+6yQjxv8AOT/+rc4DT0Sk8hVN
xKgqMifgxhbU2YPEi3uiYEsfGslswicv0dEiyNJ8+vFoDliTBMVn1SQr7Cbkyld9jkJfM4WeUdZl
5TBJMQK/MdNPiDkYDuxLjuQSNPbw3nKsRCG6Sf9jCJQwBA2MbLAS4LkkT1j2jMJTb2IAmwJQXY6P
7tduvip1RaANKYDYZuveeV9DLkDsm4Ks88Iv24hmWrN4ZT/EBNGit7t9bUrQHWCJCWuvIaYWiDCu
fKhIVKnkm4bET7KYaOGtuAZ8k9axTiH8/C0Q6qOnOlPavNdLXf2LTxxjH50gFISASfj9Dul7v4nw
LPgJkfg/LEWZ2mkbplIv9AAKEmyorR/E2DQktUhIkqpp/ZYegNQWqMR6AKsspxLQI1V/sGh1SoPE
j8mMN9img82DUQpKzPhzgVNwoPp25bMU1uS9IKqk+xoO0f3Lp7bQYM8VfKV4QOhhQkbeoKCLKhaf
DbKLbeAlBnUgkiApdI2bxAcoGe2AY9sYqDM+cyTPdiuCNumOnHzBHa7qO5o9n12B1JXqtfTc4i0b
MwQ1zf9axU1pBkvyLrKZWhU04XFxz9pdpMqyJzOHtz1idNjKesT2PO0cXAuAwg1YH23OnOg09pmW
swcddFYqUopTVR+o9Qai1daxfhXxPKQt7xFVHZmYegCq4nkLon2GkqNOFfaUKijda+7eq9Cjx3yp
47/bsgsYZyklaYsm6IC076ZHV0eFZSd2zmDKzmzCF8iVXzVgnN0IRLGWkFYUkDVB16qHzIYYsSpk
jmv9KAtkF8CaTAJtTc7ASgeImWaaFHUmf6GqX2h1vmQqBcmw8k/TJ1XrVY9mLX/hQWrxcEHxmrCs
SL7FRvSP3FrysI+2S/EANv4yKBEXXuD6JTeywNRNyifdNJIf5XQUcI2ho8YeNv9gdBoAy34Ib11Q
zJul8/IoOv7QNTtpeVnw0PPELxRyut1zFCEBdKtB4fzOrrJq+UgJRfq8kPi25Y/S3YV/fMzrXcru
qrJHQu4PHQgso3ekYy+cqpEwk02ICJVgayAvjt5Wch9ElbewU0zDQmKkZQJi8F2t9Kxh7TIi/p1n
9fnb/MBQ+WxqFbgteED/+ftXbmMlRVqjNmi4DA+2LevOW4oHXqTgqUAsx8n4+XByRKBzUMXv22/2
cdZ8V7FoTjEeoG+0v5GLbqiEbg6O8HNdWSixe13NAdxy8UQ+dGcLhZ+tTSP6+WMXSQAB5wh0tlyI
REdcZ+VoqMqvmekZ8sdQADxwP63aSYaRjgf9aYZnS9FReFs31q7hGPQ0IvgM+EwkCdBgLL5zG5Ui
1zgj6tPE/hqNDn68p6ASf+/QwCLxuLO7jD4cVfgXIhUZhlBhZDGquPzZP0xj2R5gYLivGmwI2B+N
M+VoPJWrhe27c0rcPrwU2+F4oBCUAlmDp5oPb0w4hNFr81YVIbDUuUjH8njxecziJ4W4o7qVMRv1
hIZKMImHpWeSbs+RIiYvTpyb9qXYnYFR0DAE5ykzuHgxTWsICBtTl4Yt5mZKJj/r79N4CAZhZTJU
tkoFwO5OI9mS7U1jUhMZx7Yak6KG+O8CddyvMqXRG7unOJYOKImTWsGg+5ZUj9wha81yUJLX6YaK
7SN+n+6DONMlIZAui+0oXIjodl91OW+zMk16tRFUpx78/NLyTCESgB3Ymvj2kEO16t/wlXmI9h5j
Cq/vwaynPOpUiUIvdlCJ0gWmQsCf69Q1KveJy5j7B4bS8jNYzKL+FtvrWsH+10LnGOPD2Z047RJ1
beBQNm5z3PNb3toDq66BORVSKvhSqsrDgO6uehVn2wH/0aAyDGDlDDddi6TtyOFqcOnlyiLkVnO0
pk3qJXNB2tY2weOCZIsK83/ZQnubR2fPgXps2D+p7duASOd+8+ENMZ8xUALql3eLF13+xkJU0wdq
33/Y4nP4ipjKByCbkTFNkiAUloRiV/WtNzRmOW/vbAVBmd3/8dA4tfCko7NtZYwxivDdy8ZzyCet
rQ1uIZ9TVJT7L4IEMFHNchJR2MRQgTx2d80Qjrj9TjNk/SYbKWPS4UnSPMZnSsuxFQMMj7dFyQfE
vpieh2PN4Vy1curzZ5j5ux9ckjwagLrIP8O14TMAXT+CykbjrG7hd8Kyw9QLCVgbeWRaUE8ftbFj
Hc1s676IbTktMEzT0t1NcBkdVf7V+142Sh1xvQlJREhSWxOHVDAXaJKJJe4RtoL3zIF6rFPjwRtG
BtoqiFIrZIxgYeg/2si83Dnz0f+Ajpm7K/GteJ6iJ7XiusuT2pWXrEYI1giS6S+naxX4pgh5sbuv
UV+vLY28BJWdPxzzbKSQMAcDyXeVtUiPBmV2xL13r7U1m3lzy9IoEfWDcpD3ycPZlSELiv7kmWnh
azqICbKlI9A2f3faJ4+heTPqnVcDscnn7k5Uw6Ka3MLavxaS8NHtQJX8Lg14UznflzJXqdmlNc49
RpurvSvhLgQ2a9K0Z2YQz0S5T5KlUToO0IWXZpjS4oyKrrGWUjakaC4b802SJKjqoAUx7/b1oVRF
an39qDERKTRoxJeiVIpVRWh5uPPPEAy4l1oz1ztimfElpG109HhL7qEqjdnAW5ZyPPqOPeM9P9u9
RtU6NAsNR3SfIrJ66YtKpj9sGI4eiiwWKUvw/pV1PvbQ7KUABP4ryperaTpDvTX96eg63RUjZgTU
UF1P0U5I1LFUJ7fM5rQ81z5AvB8hwjdKqU4pydyj+BGl9Xpq3PH0VtkL81P+92pKZMTE0eP/f6LO
EAc55Z9Li2baJeQh4QWXlB9HZTIonXAzroi0vuusG59Oq/OE9fxspt/kfLHJc7LMoc6oA1upO1TB
6SJtMu5nCZp7V83Plv1gN7FzSSTvFOWV+hXK0cELNQwJ7IsvyrkATiFAQJNvao3c5IMnnPJVUQIv
pkrhmJUzEasGhjoQSJuHbCb6o78LmhgTssv/GiD2GXqGX6DvzRW0QVRoYIOrxzLNHnkTmk2+zAIp
pL9BMRrS16+YAKhIhh8RYpgSGQtWsj2FWnvyTvFZ+rHnyQzxe5OVanKd5mOJrOtzIcyNK5K66RW0
pme+56EeBdvPMF6QsX8M/eQfCwO7yqnfauwfDARWqNCNCEpqLhNoiXkmxbSo/o8n0TVA0uTwKUUR
sLhI43SRD6KR4KrnEhaGvspNXrQsotf2usnRWcr0N89W559KptHiPXDlYjz6fmaLuecJj5GOY4cG
CCf5iWxPoPRTCpUnjaZfPemT2HNpWFq554kQIhOeEWAdsK0FDzWEuU/8iv/2sD6Gkl2BWWVzt/Rw
/Cm1EtDbUA97rZA53y0GzGXLjJ4AhuNsO4kFEpnQNyMIHyd+aO2e+qSnVtDx9OLWiPupOju3g8GK
daDeWedX2q6YXeV5N+wacMGrc2VGyNsIEUQpiBWJzdmRzQLkoNxCpl6EwXl3uBUox1akv1FNt1cd
wZcIzSl8c5gVsMkKCjMsqiIX9K14+33OJTkdGoSvCRTxs9TBvAGgyqzZ/coFqmZli9UBeIFTCXAA
TcTvCg626N9Q4TyYAs7L3a3PqEF+A+95QWmpcBfBZExYIgagAg79M8J/TaD/ocqsD3/SBDlTiDzy
s8aUuDf8tMrdsS4qaS8bVx2clYC5q3TPh4J55pA55FM/crnGQRDgTxKbXnE4SGbxEf0jI9GJ/e1A
bS2BSFTtRMj+yVSv9Q5m9cGwWc12SmXY9WhVdbygc06qpgN/m25vPmHZPMmgbinnsPIKtxZoWdmb
sfOT/kDyUcs/JtL0Tv5t53j/OpXlXdeUa8xmKCdSQR5TdX9OCT/Ay0TIOcytY8YyN4+oqbJNBZfp
8KUohwob9bLA2fvyq7Gl5g0kU/2dfOZQyEKAjINWG7LW87yDv4cG53rGgR6fANu+xuTaICiCaIWE
o8t3ieG0/l/IidYMbf87Z/KtD6SJfr1N5CsITDLBoEx3xWGktx7YglFnpdR2KrFwm0vlbz2aHhSE
EMeAKDH74fuHgpI87gVSbvk/ogd2HP/DnKCLQ1reRx1i8ueV5+xtVgBzXF4VWwrhu5OkHOUCUFDC
zDc9oZ3dAQwAEmF3sFPnYdf35Vp2p54XeANH/I5QVoQX03mR2RA+7KvBz7srQnSHjNsBIJJI7MQ9
rNEpSI1a4V21/D4LbahAmrGaSTEwXyHNY/ZRbwuiRl9GopDt4UrZe6iYDHGPMdGGhuFbX7oJ8ulp
+PI5tMXrQmt0l2TJTbi6uQNodbYapNdO5jrwwlrnj9gYmpomtopQwkWKwzy7DCKvW0uaI3zeJQ0a
VWCP2ra61yaEtaJ4am7tQ7sdhdZJBIQW3Gdj8oBiIjcKKqyp4BalekLdki6lc2ogDjXRBBsHdghh
lxb/YgFdn1vD7+5UVlh5+7LQmR8N2lNjn2sDYxXtLqJ52cGWWW+SXlstZ608tHBssJoGcE8wiQO+
KB4oaihkKsMG1Ze4+C0ljcNlWq3iKnzvZyJlBrzKE3ByJxqRezCdJj4zN9QOWPNBOHT/rs1Ntewj
MzKYQb+GZLKk0LTD+3zNJKj+wQJfk85g/bh/62EM4KG7BRzlZw+s/oEuImJI+pOG71CKv1aROBXO
qZoEioI+xWU20Qgc6TMYqFbIBhjyWkKPJASQcrrXKRypYbsXLM7oCLJQRcAwJUOydFh0sRD+GHzn
bn76FcU6jCpiOouJUIxaFKIOthUUPe4oqIVSE/kA0CS+uL9/RDCEF34V3efuJgrpv8zLp2C7Qnsr
p1+pByu1t43b8O8JZA/nYugLRxydTq4CNSPPiZbwvLxui/vjUgz9brlXRJYc4hS877rYv14q4fWd
uzWw9Uzy7tRiyDTiDzD0+PrpwRC12sU8BgeLDLLPA2o447eQG+9OtF9gwJgyFF6ocpgHQ+tc0fSm
HNMjAGEBYuaMFq2DLBnNYJT7tN+fIVCX4zVvEbrXTYYdj7y1Gknsi7Q51UYhhgbwRxAkwDJRvXnQ
XByCwMjTawC2IH73/lftrREu4Lh7vAn1cLimxW+kmv6cooFD6J6myC96oTrf7uAWzKwdrH3ycTKa
SDasP0wgWU24O+G/iThKKEfPzlXCJsxvYw562yWNc31sOXgYzclTgg/KRLpZpskLm23DqUCaafSS
jyKY0eUyx7Nhep7cDVXLeMfH8K8BiS9bXFlbkDzO0wMAnkw4nv5I9rXehWszUO3NiBOOi8a4+hyH
DmLPZH9uJVBJeXdc4anVXjAZaokK0A8+eorOP1OpBbLla8x7TVv4QrtNJTNDlBBuAat3z607KfcB
KC2vrDuyo+q+fMNKVdf3v7vlQ2E8qRynttarPFXf7h83lYxHA9jqLw63gzvnQpoDQG6DUFTr3peo
vgj7G38Q11M5r8HL3P1vEf+94gIK0Scs7L/wzjB1h5X0hMF3xp9YXjNgEkDH3+EJtctt3BNPirNg
QR6jeSpwB833PJGuZF20XnubRMvo4E039NJuRFB4w4+9sttLEgb1lFwjRu7U3cmNQf4D4Rc3a8ET
5sSMHN9/U4jf38k7joYL6OVeS8hPxWhRzzMiviD3GW9MlT3oSFRj/gHIrRcGU9H6AzT75o4sAfOP
ceqOXwT/YpjGIzf7zJGtFFRIC55kJU1ZomndHgMnHBgiMeR5GnWPRMtNSoisbeOLLLg5+m22OsXE
zhwhrvp3G/nUpXpLZo0TV0v6QhPxf6QWn5MJbFXlnMqEsbWdTwIucu94cGd78KRbI5gZPLOxYpYt
L88Xi3zInzxQZDHrl/4KwJ7QeNcaoXACYKgtzsUDPsPd0tWkriPY2tsMjkQO5y1hjls3rUx+DjjL
gq85Kj6XJzbrYYK+6u8TDZophH9HgwuEessKXdaLmiRlGNZS5wnk2dbkSwMf8kgaGsHjRMND/Mex
LrQZ73R93vk8vP9A3RQ1ithFAPFhO2B7Fmr2tdCuQAwc6kihlv6K0zT5wovGpjTFFQ8ejnjiodaf
ARGWtn3YhisZt4rgdNNWxNABn18RaNS2iJRn0+Q9WjdMiIvbWv67JJRxrGfYKjogs1HGXi2GdVO3
b8toBEX0SnzxFk9nNSg4XK0uWkNIyMPdRbo3G2ZR6hOYt3JQY3//B1D8+VlTcE92nCQYGvNhmaVW
UupuSvZrf6EcYpc2sQAT9bSsMOr5sQfZeyAgEjxhbjvxWTIZMZlyLjkWr4WccCitQlLcTh+u4+GD
YN7axWwS32Qc2ZPwbOG5DPCRqXtYQkajJpqeXE4YqTvnDu7BEvoNgBZFktDUJiaf+i3/OmCDtB8U
E29ZBJkhYx00/gnoQbJL/oZ1Pa0MLPDZX58y1seqrhfMza7p1gv7sG2tCRZ7K4m80mzN4dAbys7U
j+3KOiOo/i+TItPPIIU97eQc1mnelekZvUf10ZhXoAdhuL33Al4lNQV/YC6zU6yMcNHrxr0MR+ls
wH1HeZt1Q7tqty8VJFzQj6wN8ClqiN0mxUOQ8tWoXGc5yH0gXeca/BhGyLOc5xs7GTp5BAbcbpBz
76KuKf6zRi7h49nk43D2vP4dnoxP0CXai9XjjqxDlxy+iavjKkcfbqU22ThukPZsbi9Jn3VSNkS9
pokPTHnFmU7XynSm/L8OvhOsnaalFs5obc9sCpsOdTvrX4FOOsQbWJWsS7sRAFVSepi1YQV8FA/u
FmP7BsF1Khy6CTnI7XyZR4hHuBzx4G7sMxDaOCPckHXbhF8tHvhd0jUsxq2TJKXcHIeoJNYR7J+h
oExyn8UNX7HyzM+CQKdcorabaERPzHeluqPawvRvJbx8w5Swv330vd23GjL/sALAe4XILEEJ9mAM
+5CR9sw9TgNakDMIHTzIdg7nai8spl1FhtaVCf9FWyDiw20CcWwKFYOoJyyoGpvJfu8XEX3QpTpP
PPCRJ1Zh3MGBCJg0MMWJVRqOwoL/le9n00aOSZNDxBWiR1ET09kVlO2w7d+qxc0vITsUEZQ5OYG1
ohLvxv6MVWzfAe82AGYkg/iIrZYVP44/T2bmilK3pE0Xz+7eCsiQyRhaaF1FmAHE9gRoh6PI25hg
92LUnZ/psvIVoc+rPYCa43vlgGxQdQbnvrJCJzFiA0vwJTFx/dhqk/sieF6uDHk3n3zuU09Fb9/q
8YgNk5pznIQzO1BVBwcVQj8LxkdFEdU+A7yGZ8qlOxfiyY6MvRIo8yYO6K7VRz1SIU39aEMwwu7L
ifwnEH4/Or9duJZgO68/05vPQwcoMx+F84J60I/jRkLwbR9GK46zDVG2UP4WhOTo9t8sZtfwySH3
cWNZ/m7n2rjzzLUPb/MZrlj8dmklWeUp8X0W9lD9JQi8LxZKdzAmZkGNAkNbv1dhM4JpX/66dNAu
PorcKerAnTiejWBj9q/f2xBDqDMUfhDmKqTuUqzZxvk2sK2aVSvBIFUlq/akULnMwfT2tYX0QQB1
aDRrTPe09srfQ0BIBeQ0RpB3eWSO/6s1gQTSMyRx/7GbhMFYzz4aO3y1QKblRSSZmL3R5jz4sM4d
UkrbvnyTmufanNXIXM5oqZTxHCiTx8wQ7YVcnJ/jO2Hbt2ewwmEgh6JSHGcQVg5nKlDTjjdYvgin
fj3GRD5jt4pOUHB8cgjFG+UhQ3NSq0BT8CWrZZ7qSKbQw/IiDsEWKcEX5S7O/hoAoOvH+FhXs7G4
2apHoL0E4sKobfUijZAamH4PF9w8vrdOW38Srg7fXzoA5/DPEElGwvRckWqBZ6CxDMpJBWc0kG5b
A+YgAN72YrGtlbL0ujcgXgOa9tpbOu7XtmlD9V5XZqfgVgHQiOLrhPiZOZwVND8f9Eb9B3sqX3w6
Q9TMVjOicgI5WZjdx5jNAejU9y/R1wbh4x5mtAowzEti8MKLLRskZ6eggvztChiRrH9yI3rAzwDZ
48Lx84uuq4YRsuO99w0XxKkRGh6GAS+ktsfdG1TKln7OnAoSxF0vBl1PaJbgfcIESxPYaPZDy7S1
bcPWQx1yMw5kYfBGwtEYxolL2uhEE4fQdvOnrpgBqrNjltWpeRrn6KRCctB0e4dH6NvBoKh7g73+
5PV2l/79z8ajbYnHvogdpwUmbb/uXAAUPPdKbotMSJj+ypYHO9shygI8EWnZ1UKi+XdrcBUjZIue
hPtz/T6XeOLs43OkGFHCMiXbVU5DA+sR3M7DEuix9v6qmoH8l1GgAhg3Y9IXAQk72C/k1e1YoIga
Xw0mT39Yttpqjy1RAFQRvKkluitaIuqMBkrOGwH4lxHXL6db4s1dWniTczs+U3CcuWE6+eeC5oDL
/GYKGxV87nPAtpsP/69emXGqmir9gZVJxxCWs2/vmCetrraeGNSoBNdG2Rdl4EoQIsfzjS0a9N4Q
r81/oDgm8lkT9vQzV9SXcczGPuWEMMC6KZVbsiEhVILsav9F+uubheEBwBORh9RcXPvvD+KGsDnx
M6AXbrr8JOSPXDdsUR9MUf30YcZMh++MZ4t+xyMjXNQNZ6vsgvwxeNrp2kB+EIYr/Z1UMD1o+BDk
ZvKBRdxA5D7oGEDbbBTi1AImInGqFBv2+++i27lkNupTiTNiDNTaPYAPt46rttBJWosKCw8nZTrL
8ZkDOe5ZB4fDv3nK2xllPZZisq6joeWCNXcg3cfHWonLYAz7O23zx8WOtnLUye3RllSGZNBb9Jzn
pvb7XEFUd3r5jrpTBhhHGtY+M7zSZGRWIOpGp0v7kOgT/+NVa4HaL9w3vSIutqzi8QnM/3z3Xspw
IZVkyCsQnbFXr+eOkiPet3Qaw+KQW+dC6lcCSdPNzZnsw6r/4neVX1KPU0cQ0oHOegjo4oYxrWF6
plm6+BY59+fRv8xtFdYZ5+UNntQvX5Hpgrf5EJ/1JH+HPSKTu75m0HDmoM8D7v1LkaQoBj4T7OVs
Il98BNBBpDkAbmFKvzAUkOXyVmYhMNM/VJ2OjWEq0bFRbbV0aZCP52bvi/B9p6zJg5S5/5NYiUSu
poj71lKetDw/2UciajTIhYgvMr/GeNnfvIcCVhyX78kHLIQcsfdMYU3jihAtcHzMVvROcdJp2XIm
anOcaYLChbM3W0FX7Fhik6BoJaF1o10HrYlkgL/fL2lfgRtN96hQhJtKMIYqKGSjRFo5tVzOriaa
qqyaSZc15lNa/GBM6qZQ1ntNcsnuqPvC9on3B5wX027F6qcK0M/mNcSjAw7YRrHl+sGp4C6g7xBG
ZDfc0s6UpLpSD84cBw5YZBytk7KtGXGZBaOqfKIqfMwBXnPFlIGTyTP2DA3+7UY5gBHeCnUWOBcY
p4DjEXFCyy1vEP0chmQmMDudu6SKkzGUDjP3aujp59BVH67CKd70yRX4nPTuCByIKSo/ahXJgksl
nCxi+lnzuys2+evNkhwLEXwyx5NY4H/SojXiGpdUN6y15qReI+ABwPDJui7Wdarb5Y8LaQznCKmD
LM/G10KeRi1uuHMU+ALLSSg4t2tOK648yERMx3TPNIGdh5G60cNLx/YoH73J+6f9rwNaze+Xu+F4
UPCreuAxZshQVQAclrsXG+qlrcbQ9Z0X7cI3ZKltwSRNbwFBRcFM2Woh2HlO1dEoxggwJIpxo1Tn
qHN9REcJFHFesxbp2eR3hto8G0XCWtCT4mqgrxf0wWYagIQ+aH/ZZLSwS1QFwj+ckejZAQhMNSI/
r4m4VGTy1A0PQTr2rzwSg8Cmz2QnAOuJyEet9RgvLGXLQBM9sZZWd+gYCGvqMZylRp4hHJQoiJtr
Al3aN0aMlCpTazAtvkc+O6EPr2yyH7DbHAHgyu/mVs1NaYDbvKQSNND6c4NFORHL1QLdo44F1Jtv
UiGY9DLMNgJvriJYaEG0myzdYep1QfiYG5dKcBRXpjUwVUM9q5/MEEv68IJrUBhGawKpPZ6EiW2v
XTKwGhYDFaNLmda6yYwgdFD6In8raS+vC4Y0rd69j1H5EIShxh82Dzv+aTyEe1Xyy8czjoOMMC8/
v4OdCqUJq5C5oDV+VdgMShXMNXrEvIgrsNj31OU7/0wF3NTAYQhIT3hOTJ0DlP9gdjqTTufsqsiq
nA2kpqs9nNUo3tVzd1LBefibMC3VAGALmYwvjcGquz5b3NHBSmaB55rTH4BfBCNpZQyIKPqTR9xx
h3E4zbXsREUBfnoMYk/B3gDkvEMwAKjFuBt9aorsgc0NInj7GxDR68HlI5sUZe62xrU4Xs480xnm
IJh6J+N3X0+SX4K917VoHEmgrVOJuR9lipfltf0tC1s1i2oU6arZtznQpksSptxi2wtojKfD+60z
4OIoN4sNCQ/Y5nJ+dxbfpxpX5bWLXMNxyZx4Vo5RyLs7Dxqw3yQcp3vWFtvd3rqvjXPVwWgM1Ce5
CmpI5X/MGYHFEBnxJ/lt6602hjd4QtIoQRcC6gvgfK+f7/vdFuNT1dWUBy/pFfBu0v+4AtwchUkL
b8MK8UMMKloCaTjMnDN+tuc305wdrAaj3FMzlbxf5xmsy5tL+/WJ2rp/PDm940xOGu370T7UVrGu
sfNQitAt6PdQKNMO55yq/0cHpr2IrWc9wb+lrVQIFBJvrbx51rMzU+ZjdSU7Lhu12DJG66qyyq3+
vTFr0b/hOrX4qzFE2G4WGCIgA4w4qb3aBfXNVMGKokDFMRW4fR3BBjZcZj8Bk8UI7Y/eMGJ0R2HC
pLMoD8LJmcWYrCbisHUh1JmWlGceSuf4igHT6fkHvmWQGuehw0VJ8cV51inHUfoj/7gCZosFTXcl
2pvBxFln9UO+3lfr0BL3IqXotGNwl86MP+gUAe2tHu5jCQ12QsBy7TO5B5wZA3NI2nl+xodS6yaD
QE4ADYp4qu+ZDHDuYxhScaAo71vaUieCpZFpKCkEGUvtj5ccsmLF+11JX6QPSTsj5K0x++7mX/sa
ne9z/ZJQ00nVD6uETfSgvJZXJrzSMUL48dcSiK/QfK4ACDPKkD9Q3fu29LbnVogPzP1me4ovL5QZ
OuynMR6GL/rq1bowY2GxMTKXwn8ubMVYYIaGi2upoP1slIt8oH1dWaaGzmy1rFxwug5TGnVpgHeJ
RYec828ud7BHD/Y5UXt7tqGzFaCXMpbAmmwQjlPIIs6UJYRZztgJWs1n95Zo/WvsVm4JkfDPRxpY
dwCSg/tAjZkD14OJ9ZkXcrr+bYAOFLMtHL81BcTcZnk9pIdZ0G1OsSa1pmIe2oXlyJeHGlUQ6FOs
PojA1OCedKXMgPxp5a9TnRCc00Ku/7GGx0cBoCOz1yQYA5hWULCXf0YvlkGOm6YWdeqGirtTZvlL
JiyWY9PydWK4AcnlWQWWCnc4+r/FVc6F+2/eMSj5mPH67NlGuZgM1VxBTfV77ijrU1hTvTG7OYFG
u0lGFnooRj2kjjM4b5cMAPhMSPeA37rI6VYm5s77dhe74xWxsURlDriSraxPiB5BrTX7dnP3Rz07
bHGKPYxW8YrrApc6e17Z7lxAZfhRYJ8GtxORbyPwkIw0PBG5MqL6LRkSF6jM8Z3lfwGiD31RrLL5
UFAa+A0MXrwQGdXhmQ0VDVk2iseVBplQkX+LFhgbbfkyKlLM2177JkFHIe2KlIygLn5XapBQQbcn
P+np8E7v21kmOjVGB52Vn2gQ/jxe4fmzzVMtDxHctnrUppNzWbMoCcFMvzWE7Zjhj9UmLRi/d0AV
vGm5aAyJ0sY0v8zprYz1B/XOSXvNQYuCFdlFKsnSAKaXhH29OaLRT+eHhtYBtVdAypZ28bxcmZUO
svjMP5omG2zqnCTsQ0/+MQXMlJ0MMwQbDvLBQnFZL5mTtpvDGo3ZWCqAPOjwDQe5HU6WyvMyEJrn
7J9nJh3/xKu4QrhDJWxsIwNcgbiX6kxXYyD6Zw4W45w6Z0WTzuOys/aG+G0wYIzYrdbC9yQP1SnL
kDWDs/FjfzNUxNwrSJBoIbbPkcG2z8IBFtnxfGstGSe+GBD5K3AZTeqofjfSEE68D2VTT6m4yV8U
A9Ut0mSt1HCSgekc0Rqk/klUKAWoZHnDm2+jxNc9ptSL28qhzlMbxMVa12r3Ka89/1ZuzMxzr3/s
wX7QmaEErgbEoZhz64oYhsULUqXj1OyAMT+J4tJOIYS4r/bPv71meNBvsvSoMHY4Cds6w/9Ur4Qn
glmF25Os6SzqbsUYPc+IdYX2Y6VsZ2JRds+EgpbM/e0jDAQuy+3GIXejfni4RflZ5MfjCnl1nrSr
KwxR6jrV5RABP8Dm3LUNR5v4D7oQcbpLEWq1ogXVq9ducEU8wvLOrcR0S92xcDu7PkL3/Ic/CIWp
9wn7UQ1Dw7JCHQQKVzLCmuePyOsHn7QIWkzvAaWwVY1z/HfOQUq3pMOjDe27djNCCPCxNrnuC+Mz
wuaHKkEWket8rQqvW9iXL1E9AP67MVh3SC/Ofk+ClzgnGerlsWP2tuWiNx9S/rjATGp38C+Z7bJi
hy42JArqu0YpLOB/fKZT+Cz4My+u/Y7GtkPGRBiZ5wpHa3bKm8SjQ331jMLJk9z0/dKuqUbcukHy
HnPhMr7flpragfxeLk1/8Xt2Ll/dUAv5WM00hKfnCHXohKehAhcge8sGB1GVnleYvRu5w+kIWGyg
H4o+pK2Pi+HbvUWtah2TUhQ0Blggoch+LeKTdeyR2IBKUqmRdx7WCylrLxsj945ZPttD/mzjmfyY
UpFuIRchJjMb6hUd+LB1OAcFnx5jbAEDsg5vQEqM46ze5aPB3dERvMRcPeUVqw4cNTZy7bWFnaEO
QFcO8PmjZfKu9Zbr1mhRr7DM9eaiZ+UQU8VmO+jQxIkVoI5g/uRJ7Eh0wly2LILtOezvXszrWE/9
w7sl+UXkCa67m+2vxkyWzV8UvUhh8SJF0BkGJCbA+7vDmvTy55tcBJH8qZtW/Ky6ui4jZChSdWwP
fkXAYY0c5oP84OaYiv8GrKgc8t3YyITW9YLQnTbJ/pXzewPpmAlaTDT1O4XkK3Kt5qgrR+gUNxtv
Lf3kVuR9ZFpYmed1eGrePdQkEty5S73cMvr9Hf0hEwqXUteUdOo9V56FR26xKNzPOgrPlFhM9LgD
ru2CWxePJmHCpr4aYYsZVG83o4eR5Xu18F9+sd/29MZUh6cFXX+nPeTxqGxnEmR9eToPEHZxzkcf
COdL7Hv3GsNXzpz+QusUB98wkx3TvkmNvzrZnfa1jb3q7ZtDT4hW8JkYf+AheNB69V1gcTr64/km
r+a4Cwt8VqBvX+qO/1ftfB6zbDLm6Q1fTtCkmge3FiQHTKgJmOgrD0YrhYcqh0g5JNOh68tuWGgp
aashn2pl/wy/5Zp+evlJ2KxxEa+UaibxLV5ZAcDsxiw87maV4IQSKIszpS204GKnaMqdA+aBpBdx
uxUdp08n2PdvBhA23RSs7JiLAyyNX2WStf0iweDjVhjesaN8VTJwwkDQUv47JhzYtTmVxNUSP3G+
2d+5mKoX2toAiYD9/PjEY3T0ieyU25UwFyvkkpAT4t9CvjVbzS0PEW1MptU2SMus++QV6fAzFDW1
m5vUYFAlMhRMPW3DzTQrRykGhgI5fTtrB/B4ElsIuVhXd9O583r+B8ffeqfjMXkFkKUK7z6P50uP
EV8TxaTHLVaD17c22dSKUqmWXH4TpNZ2evsqcdqA5dfEkv9fvbmtnhFHhfqWlTbn0tsxGVe9iF1l
0SwqMOyh1NlAT1njVLdPIK7ggFqO1ZgJXLY7RpOe8FXL4vW8Bt+fNAvuEKeJon9DoMf1aFjFzJ0e
zBlHj/Q1T8c9cdj0LGquF0cOsn9GMO4GFOHM49HsGQjmpR66S1Kd90T3MSI/BqBhk3WFoF9Bknz3
U6pP8myBr+WC+Phov0pdpaRxtVum9xkxag0BRjH+hhVeW6QlSd7lx05GQ95QZjwhyDJfGVCYg3Ca
OSpI4c9Mc235aRw41tbMZapHhp5sK+qIu9acKpXrD63i7wz1miFgnGVNV0A1Y/o3X+DCe4F2tj6V
/4f7y8818sAwpxQ5jRnzJTtOaKrbOYlZ8zrtJruEWnGPI9hUu2SLd+RN60daXC19+DMpxaoAVmk+
szE3jDM2I/JQ0yJnPVDk5CBcSoRlE+srmWf3+JOHntt32sbk3OmwTk601CZ5BvF68Ln98WleX7FB
FU4UvTVb0XPQDXjXC2nOiQxJbd0wZxUxR++rP+piZsuMpnD3mtmYT5A3zpAHGt4I14f7dfwxv6Zo
k6nP50cTSMzQkdtWEUTnXr0LKon0yzmYFaK9hn98Qo86Se+l/IJ0IK8lfxMmPNeO1C7nYJXlkZSy
yu/Gn3qsvBHBYnKA6apMPblSsoCXeSxjD2jsNigOegwWQlv/mobedw1+I+mXQiKfOLDAzTxGGOiA
WMWxLj4EYtjKAkIFh2x9OUtPjU06nRGiXU0QzuhL8QmeMbfcO16Rt7lMYQtpKRozAvaHdY76Z8hf
bgHEY+uU02By0fY1traDFqijckbfPtYn1/VN8YVtcU8fpAdmUAd2FbSFQmEeywNSYswLYCUf4MU9
oDoIPGOkr0mPPK8GHi8J9WhtvG51SOU5xlbW/qByaodRii+OkYVYnnPotGeN+59UogiI+f7n15Qh
GqDezjVnCXPFQmS6kJmLIALp+FoxiEbD/JHfEbGzchMdy7+wE7al+lRXrLfnkufb8JeuWiI5jNsl
zZLllQwpunrD7VeKkOLb0RF9aOfksSnVQ8uBifJ13lrcOrpXJuOPAwISjiEEtoba9sCpw3UBURp1
24AsVXbRcnrG3/sC/fQmlCO+hLJJk3+1TaFFQxsFe87a+/tsC8ec1sHmZR9+zE1ezDvxvrNIC8Lb
iwj1y6US2YsaMt7bb2AqT1xD6Q7Kq2eCVd2dZeyc30OEhQHAwpIcezQQGqthtNYH4uO3IeTDU8w0
16LFSzU1R+JKSd7P1mV1lGyXiFOIsDCIypf5ZtNreLdBcr5qfQjEFUgBRB674hs2CU+/zMXiNfy+
/tIEg4I80ezzNA1WphXAFT56P3CzlonUufRpR4a5aeAyB6kGhl68K8MOvQt6v95+wdOtcY1hbFAe
PIXYi6bwE0YtoXuoqBqMGLRsv0xDykJiGrpdSWo0zkib7oJXva8bZF+sav+0Rw2/FB3dgreOu3Nl
S+NoBNikOIQzvA5NGKvjCJMgElz9It3gYk+dTZzTMnRypcT4SKf46s0Jt1uUEFn/9o8hR5IGAnnO
b27UJXvK8NPIZG5/vKKRJ9Vw8bn4UV3/NYUWbZNv0kYrtP6xpfsk8bF9OO9iCyJT7agT6jMpRHhx
73Ce8KJ8V03i07ZsKsRwNb2+QpLOnr71304Rgr0RfHZXV+a8YjsC0m9aUmDmFYOHGvLQWC1Szx7b
J1EjoKASlf/FU63L3Nb513dY75Kd29TnEl0iYGDt+2nwZ8CxYrXkEJ2QW3w6CTyF/YUczCfRlPN1
1i7nYla0DY+CBWBx5p8uwtppVIHQePVerSHKef1ZPtaavrKPAFfZGtOCRgu7WglvEZBiD554wH/Q
jkrTQNfb79KeNlt05GcPvqW+4/uRt4CUEVqRxHXzhYYPzbF2TqlQdJI5pd1EbPvS35sP2EmJxPxM
zTll6mCupt/RpkILmcgh/cZOVXmQ6GrO1+M03NOsmVakLiY0U8nwaUkPcHG12fw2OAhJ8pFlpPOl
IRhzsCdWLqKMastCm2UTYyYipx+B8MHbhhG7LedRvgQFzHFwCIfJ14YZ+ogDdv8bJcN56bvjIKGm
d9oAoj5lDswbCgMb75KJQCu4bF2H5FVvEDUramPgeidB7zZU/fiuFE7toUH8SIC/0fXhRLJ7Yxad
aB3trF/1GjcfXbHE2x0JnwzpWGtFEkakJsBP2IR6bi+Azex5f0o0RrVHqNeKzebaQ1jnCQ7rji/J
qhKGmiZxqyyRgmf0WPMRptHPu/Cpz0CjhY2RFS9rWp3sdLxbnVzOnUYlNERdM7cd+vDfccj099vX
itCV6llzcdr4FYoexI81VnEMtroUqJvOazpDp9H1Yczq8TJI19hzay6C3kocSGLLgGHByynlEqxm
vQZsR+LEnyFURXViEQaRHteXs6g+UW3DpLw0Vpc6zgM7GRd6Y5OGwUtIVZdGv0ZqMqELNtLclw76
th1LxWRj+6JZA3Svv1hgfwNgcWRV4+SKyvpGJGBZNKh3g8f9JN36leO4G7rn2rl4eRzU5Ssf0UZY
WB8g6PW2/EpPfq00bAa5hexaYsjszqgpt7HRK3xNY2+g3s7H4pmtHLi4g2qvTZZGnET+CZ4Q+BkV
v4WB5RflqNysQg5WakBooDavZil6dW48LmaHbMopsUg/SE8DERRg52b1aTd2kKFBBmpRFcwxI5dP
M0Qi2PhMCP935eTI4xCTDiXGwkPFs+1e+Xn5WvTu/0FhpHl+YI1JCVPdh2GEifs3/4cdZJ9ntmqg
QOLKluIRuTsjXnYTLBZuC678d/5ELQQ9v7oU2UNjPSXqF+aLXZEw9rQuf6yo5EDJsaQioVyWehC7
ErsUgG37Oy7dI9X5z/Impik5nEUB+3sT0nzB3xA3oK8G11+t4Qq7DbjOAiAVPy/wLSxNuUlt6hEw
ijNlZPvk/dEBP3W8tJ53yEnbynR8jhWzcbyZZlR+TrhvXqhdI8SKdleNqEunO8e/l0L+zM1EXKWo
Zquy8e3aO3yI2313swczCL7QuFEnoeedZsLOEQUHGSirZdFKnIKEc0haM/FC1k4u/hIkAVd0RY0U
TMhQyBNEBUuQvoHsbCswZ6Tojs2jJeDUYfpVr6L4KwMVQN1HuXa0So0g89Q4vw6b3ts6CmQBBJz1
DMLqAAv98S9K/1EMHfzSoNDWhT/Z27yEgoWeUxpSCN7700mmqKF+kDY0Y1sTrFY6VPHFtb/6iJmk
nnJZL1HK1tQAfDs0T6UWDsstI/W8skusZHchuxrMCQpH5BTxxuly4DYE6AOF8rwwMCyOkbJ9bokJ
P+DLMhqq461KYRzPpdNz+pBpIxSZNf3eyxtdrwK3JUWQ5DJpZ+/CrIRh99fXZYmr1cLtkF0DFVuX
L4RS0Xnt9SnXi8uXLcIt7LsrGfvz8JOb1N2IDVrZjc1bwpAfcuMXS2bjCQQyemOV0Cv1gfbF6Tqz
Q6JgeFcvmcpK0o6Gv9iT5UaFdBoc3kPiDRrw7TZzlQFWNBLdZMCo4Yt5Rev6+OQh80cWJPBcon4v
3sDiFYyXwjDb46wQBGLlP8nQReiYWU4Lhm2n3uDBmQ+qLH63cUGqlXw/XcohFwk3a5/xOYRp25I1
P4vuR0g97jSrt0O3q6XEG5qGIQ4swmJ+ZKIbMx4qPcDMr/bh7K7QQMdfr1ACgUqOVgVtZP2wX9JY
BAvfgdM6xs4tAxS5gLN32M9iScNJyRirXYz67nRnCV51PPOmTrYLhNMMpGmuh479WskhjKvMYeSV
rTwmgUiPwMJSmHGRr90u4EnYiSOCtfXWkIT2xHCUkgYs64mqtFJtVsITD0RhNo9ViAqxGJ/mjUE/
8kVnzpszVzAzXuW3ziLdoC5EvqDJQHKcNbbLqP38poJc8RVmDZS636mg8FT6rDaKriRVBTaycui6
zmLRD8zCHaCCeb/Jjd/ibF9RbR5eBoVQKbvGQP9kkYtAKUWly8ky2q2Ki93r8DEkO/GhfmV/Mhnm
VRmzhYjwA/ZokBbSi9pbGdxI3yD2zLEeojiU7Yja4CRhQwAAOR4iL74OBzxV/wXi2wK1IZG8uGN5
WwVibij5sb21XdAjF7DZcL2nwIvBsxSoXhdQe1E3jE8gceZCHekZkEJK1xUFP1eZdV5AER4DUb7n
Bz9UGWBogmThAaIOezOuX3kEg8W7PIyA/Sbs9crupBsjwEC+nSSpUaat8IctgDmB3kaxy7qKf2KL
iK6KI5+Z6KSC26J6gdM8YQF3cxXB1Mc9j5oyfBsTxBkkql6ya4ZYWSPTAV2ZuF0DZcbLdN2a2tI5
kmLHDjGB9EW8PdgSuf21PyBB9ojtagPlFoxbIhA/yBYmTH40GAa4j56sx7v6DftN0m2356C1FmSA
8Pg5YpX0jyZq3TL0bQt5+5R8GSRKufO7n1PGkS7FvTv4QjFXCSq2s8nMTs4cuREdXou4pwIuqPcx
WeFnyR43gmBVkfV6lI6v72tc+fsDtZeemInFNCDRmE74AasqhOeCBe9IYYq6dT+sE7W2YlfZs2fj
Zk5bOwWsaYcKVaTcpaY5VCfwV0I7iOWnRx+O3qbSZk6FEr8l2qlH6SJFOER8JDa1CSDvjLCDiW0d
LNuvL6foFRYzGMnbm3dOWIjfCDLqD9Aj/kOs4xaIpUJGAobgNnM9S54J6kQRr+gqGyL8YwtNd55J
9bhMTHNESfiCfrcmGCEHO2YPlmeZ8XFBTPdS67VjyH41gSY+EeFsW0Dz4QAecrtfvK+Gyq5KdpPm
YJzaDVd6goPpMEu13xalV9BS5Ry5UcJUjuOlBBERCaC4HCE13/Jdlp5EfUi9njF7XMCWX1OJsFs6
eb3WHzXIYsgp+7vi6plOkYAHWFsZLl22KPGyoigjMgYvyhhHTOh6ovfgkNeFQktILy7OoSVp58I5
ag1IQ1VBXh1XZlIPsaWahO/mM5Gku+e/l3ryuOu7wftDkzYg1zfy4TCv7DRpBN7qh/CIkMB/yIPc
cZLw+G+ClZDZZc7SEGkXe+Rx3kjSAQcUtdplrzxahwTbULWTv10p9GbTcxGqBIdlo8Nfrkr97xrh
J+yPKb1B/IvpDfdnejsEmIg+RSxjJY5GG5Prz/QaWeg9d5D7RvGYAQwSbDRssItcKzQBT8HEThs0
mUhIXm2i8g/F6jnXK6wcrwYzNVQcQ23AmpbwZnvj1CbnaU5AT9iDqgxaueynwOxzqrttvRoxNwwC
/Pzrirq1Lk6RAAb/6wI3gDa8GdisCoZsIosdJN5Lh/R5aPiVVG2cLrxw14CvY3baAu4aR95kJQPm
AMfybnhzdVQjpnl1sZ39lggG6a+lzMrhfdUslkeStT4tIg1c9HHwuOwKFr4/Y11GhXyZqjNPzO+s
Ktb9ZZ4X5P353NlwwTXJnzlYIIFlGvHjelUYZdL3CcNzCQUuNpNrusEjksp3h3x9g/Htj9oXkOAY
IWvODCqJKG21Gjswn40SPJMUM51FEYG3ikYY8VmZJe+Iu65LGrc8kibUtNxmGsmD2Y/hFh1rScid
CrxJ6/nQHqnHtCm2mhKu5oDmmAMEXosXxkW7b0h65gngmzAHe8GsuyvqTqcRPYx/LE0lo0OQSLIW
jJVhHH4tEzOcbDHsWfzYtF76S+S6YD0QEFrjlwnOpxlqKadrGyMTvYcTGh0+mmnilCg2mq2SIyE3
Qp/Qhd5K+OeJvL7HHjf4ExWdxD2mAub4mspC3bDC5YStetUdW7AGZFb5d2bz5ZDNbyBXkz0Hp1Ll
o9WSYSQnkwCzeGZ0wvyav30Nvf2AWUg1DFrN3WmvooBP4E7g+pbBOBXe7362h7CzzQ8XVUDcZAnS
+Ix/7ORPfEsBWIlqp0hBbgcevhNE/64s6J7QWK0+Uy7vRklq4wrIG9VgV49rUV8f4hLKC6GCdb4t
t0UqxtMHQ9UwN02aabd1RFuPTd/ekjGZTs2yDUoAjCqYq9pDI7UuZ8YT2H/rn6p1Wu9MwM/eGFov
pUEK7BNxfKGgE9BQm/OTYVwty5KS9SYEeB5uEoNXiH4sbljC33b6ARwDKboEyT23FJYSwUFTgYp/
Hn7lYBUxg4KfdsNZ1KaOki5eDhTGhrNq2OwngCvEYYLeid141kJKZNr4icqGb/B5OQ58VdzsEDDW
aXsy0j2VLK0weK21DdtVy88JXFPO/8ZMB79hxMZowBexI8tOn7qBNXWcILE0Dt+GlcsEWtqLb3X4
yEQZGEE3eyiwo+3xAIkw8QFhbpjQ6fBdrJ90V2f4lMdzKgrABx/WshE5+ZAjG0/v6Bz+6qh/0t5H
LYA1/IVEAS98aiIBvUbO47r0LCQYKlLYHkqoRS9Co6e0YPqJAo54ugWFSEVDoxMuxNQtar20Qu+q
Z7FirTuAA2UkTlPzqU6cx847+Q5nJUP/J3sNuRznTSzxv2kpvs1j2y/kTTF3el3VgZ8JFRvvewTT
tnpk3dTdoWPUsYBC1em3qIJzjJ0RbUFU6OcuCqgWg6y7aFJzznqanxWudIzdwPpv2hotaX0GQO9x
usCz3AZi5Ar9tkqzj5Qt7f9MQ2O5gA8AGjFmTzAtv0UQ71lDvASymn/YwtgjkXDRK3JlQIwwUkp+
3iqyEhicZDchfoFtj/2MMgCUqBG/sg/3eeXFFZGf7ymI7SS9stJ4T9uF7U2eBmOG3tbujKIL/oa/
eWII6has27foUppHhtqGh2z8qF0335sNEJXeEyIBVGMlkaSmNrzadoODQ9xd/NslrxO1MohFOAvu
Vm0RYXOifXafgxmikNKZGwY421j21/4Yb5sxhlWHAMXyolHQerHvptamS145PdwTow+lk8SiwopH
XX6zvm5lzehKAmyx9Tiz6TvbmDup4ytdu8nZJiLykgyofGytayOJ5yWlLMsjvHfvWBEDY17izNmI
dB2cZrrjuoMIrm/THIWhBq96Ok5F35yLXz5KDuPXV+DK2OK9UfTdsmT7OrOfegqIXeUrrAexFJUS
vNqO6nqAX5Jnfr6Fl4pr4tVz2/UMaQDLawBcijoPsHvkRzrdsShfDdNzOP77WqjNdFeop3rotHf4
82wzpOkAm9UcygwIO6Y34EYe/Lw8KqWO5MN51vQiEuqpWSPzrS0Ii3A1q8tyy0YhT1l7xoePp3Wq
CGs7YOLhGv7vNhTbTpmCuUEwYO60wJsq/ibTXieoyX3IzTkJZi6fdTbr/WFt8gCIi2GlVn+gkSC8
55vXRw48cxWrBoCDq8O+EO4BWKkn/1QLq4uGeijeSZ1bcFOkd3IrRVHubbkA9ima+CXgGbidl/hc
9KEX5sxyigfaOLIwAOZgNVSmQ7OOWsxW7GtUd13/lE8S02a/YSAKrQm0f2dkEcZUjm/b+E062oFM
4ouH68i58xO0yABZNfUU+Wipw9HY9kLltAmqTRrmZfzZZxWcLiDT5qFsERNLGJxlpFiqMkAmggay
56ygHTnGovxDq2EV2U5dzHGa0kDbiAWOOd2TU9HKWVNqXoXaZpZutg8Q7Km6JPYnzEFhw5p15YRT
Gmjprr2+QaGcnXXI2141Q2wEUavSg5F8bkgZYhZO6eb+IfXrHyJC65oY3fsqMiStOtVYf4ai3xN+
ZcAXPvDKxp/gV6NUhP2VagNEKvO8Boi0tW1ibgabSCyenQ1JszIPVKklAtMo5di8UKfYnudrbgk2
ynC+5Xf2m5MB0nPn+sf9qK5PZL5Lc8Sl174nGat6U4zoydZO7kjo/xNlD/tYtCcX0lMn4lAwkCEU
qxkJaZu8/4QZUegeet7HwZ08ZuZY1S2HO8TluFncZwocLqbKZz0LxmNRmZ0zVmpitMtuZLulKcHB
/Ugnb3IOjjHuID9QF5XGh/KiT3c5IZjeqeu32j1sIfKmB6Pd/0+pRGObDqeLcbyo7rxgLtNNWC6T
cUZcMSgfdVFe8MDootjzgCHTJ/DM5w6kF23FHkqsKS/KgNCnJcCb0w7zIe80kmwq+ug46BGX2dHU
SLAkdtcAeGQOul0C9U1D8+izuTmdf7fgm22QgtSFr4oO0DFVlplt4Hgqy/HJjF4PW3UBe6ar6oA+
qjJ+wi5sVj1MfBmTH1Z7M2lCrBmoziZ3Pbgle4uGqaJzVsGbKpDRsJ5DwB3uAlIGzOeuyMOnnvn+
0oO7XZQ0akdgALbO/1AnjWdWWdRvDAFMKLHH/vqIr5xcBuYpwBgmgFiWPq/cAyyDU87dxZnHqPOG
ynFBPIOlU9wFvtzDt3AjLRiNl2reaTw/BisobxcpGKCKhZdYABGiVR6JHsNRbmb1ZaxwyzUetOhh
rKSujN6mKo1V7kgisnqvdpCRe0hFBdDyixmFbXSCR1la/l60E4JfJ3LZxowkzjMLHtFj2mCMnAIQ
7K19v8wwjcfPYBsnabhwnNJLQBHiWqjK/V6JTWNGCLNEs2V08b/VPkOGY9OZwOH5UKbaH3R8qlJH
83Dt9SlqzLSrdTxIetLZfr35rlLWsoxBYoCU1tJ/yqtxk21DbtEBE59/IiQAjvCPFU+owIL9NtGq
LNR6OIs+wNV6M4L+irrG69xn95oKvv4LWvQlgPZDlp0ZSTUuwzyfYKP+5N+4q1dfEljOuAAGmti5
JYpw3pG4mGVAmf93zV/7EZ3eOEV0IKL2/5ZQmOAiD6Sxgo0mlPZ2lRMwPLLYY7ZR35r4Kq4oLgr0
FzDfY3cPbHshUFjVQai4lA8+xaCjCLqjLJD6fMqyhx6moEog/sSfQSgRAwXnb8bjzqxjAylAUD+B
/qbK9n6j+nMzhpWzHrBVaCPV9vBIanSjnDCbFreoVFmU8MD4yz8/bcu/3CJbyBwppuhQgHCXIOWd
HMqI+V5/CgF92L8rQlMcE214F2LZc2iOSPuFYckfQP2B7NayVW0SEKJV+dVeocIrs88tgEZDePVn
WtSGJKjQkY6nji8rS08YMxOqOpkD8YuhK8IWG00LuyhZ3K5G8NCvCQUMGbzGdxNmbL/66WtGojj5
g+9EIMpUCm0GXXuB6vlEc7RRLXr90HcJpDzIh64jyfxmDtjPtfIX90RKI/D8CCgZEYaiXV8QmU0K
+ovDJ9q+G9NW7v+wkhhgvkMaCyZ5dLpjvQWbq92DE9iL4esOSU384ZHlIIcOUSWItFsVWWS/Ofzq
2LsmiYxHKItfw95r29BxOlNLEBnmDwKmeOIRUiHXBhWuLcRsSUqddvTsnIr44TvhaNmhYLP9Zc//
gkaFFOgpy8DjC4szPJ1KA9J7szouMgtrMAkhz0HXLfp6UsNpGrzw1q735fITDgZcaH2M9vibO2XK
RyWqE/ACP3/T/LjjDe0y7OE+q42ece5gxFe65CtOe1ytK5xjkQiZ1XiZobssvSm84X41jYMrHXKw
BvJhd8CgHBIUWcdh1SbuD9ZeStTHy47Pp5rodKvS57COmDq4y0YpJzNjrVPBupUjPqcatjrLYKav
LSDuts7bTU5HRid1qSyHqo45morGroRleZewzGSSxOyQ9ij477A6lI9PHu6eL3KTjnylSn4sXecS
l9ec/SuQXL06oauTD7MRjwbBvnF+nKMdj/gmr80cu84iNV5LiRsT9WKunA0TA21gqkfc4RSddcwQ
NATR0I8XUAFmsnq2E/HETb+eupTmHRFdIweirQEeiPNEeLdedmFIdCUBCkVNaQ9X0UncUE5nSi3a
jdDncktcOqyjMTaB9JSa2Tebah3ZQ6Nv9iw3eccRZirvFL3yfQFe+/k+d+utAfnrCsTDDoTfAe6F
Ypxjv7AtT5lO81+krs6NnnjRgGZVCOatKMK8QL9aPGnTR4pkQuZ2LPwPrGxexg/gXMmfia3i8Jpk
oWm5Gy2Wn189XMdJ0fCMoHy5ttCuChRQ3ZP/9ez6IifP7XP5vXiqjQl68xySCSr+oTWLJoHP62A1
tkni8gTUQoKyPNgtEeCyueuiN0FS126AcvnMvwJwtedUvNOwG/ub4axlylfeJr0hshQjiqwOlz5D
BwLoExbw8Fc/ocALY4yeTHmNHRczEhUI81OG2m1w8QqLkKLsyjpul4Anfd4cn0tT87UzJMY+3x/w
w9mekIOQrvndpd4KokHJHLsiDniCEjUKdup+HztDzveKZ2lA6Cxsyz5hqKqIguWArSrmm3/218/h
2Igkt8nVciMwPmCFTNYQpDaxMoU625v0+88ZasVuZM9rKfajqoInwk1WR8/y5gccw++U/4v0aHDy
JpW9Zzi6m/yY6FtfTwT3p/+zbFBkRg6h4r+d2o5b4R1lOD9v4A1D9gnXEIKt2MAIhk+qxBGrVwex
cYCOCGlPG7N4ckQMmqY8ET4h0BE+OFRv98AXrWAvDN8Qol2HJvtxkNRiJpqsCcGZ+Ma8EE0IQ38J
8IwxaS9TJ353tjkRNrXG9WfXkDejSsdT2lYlGX3NIyL3CKn4FGrP0fD4guvGX0lu7Ozzz3smasu0
mkRQHtQtbduGVOwuAN4k8k7VvJMHI96QAZY1kvX/UJwNq6A/4l1oB3gwbsi4xlIOJsFKoOG5Zf78
EXARstNR+tGyNYIzKnf/zJnP23tKHK8nTEPcHlTLy2dfYAdZ3SDQv9qV+Bg+zblQo0vg1TGrD/1m
pt0/kuFt0UqheZkchV4GcP5kInehn2wykcOt6AiuUsdwBW8FguKBgl7uE7IixbTC8oIm/PBtG9EE
e/KzD4B2WIk3uCfEEe/mWQQe9cGSqg65EvD3Vcw8jCu2VCBULUWd4mz7Ym3O+j+zqXI67pceFvyO
Lo5tmtXSY2hGS9B3etJmsOgAtLo5V/3kYhgSMBpnsgIkIcfpzawSKTvEAyZFHXqd0dS7c342DU7b
rDD/OBaJ7PZddHORZYq4Pyt6t0YTKHvukEbrVVn6lbF3e/ZQdtCeF0Eeg8ShPfjytqL+dUA+Wy9S
NbtlORWx5PUHxhWkUCX//Bteq/RfnDTaO2zTfdxjRKB9uySWCaLSAezRhJBn83DCT75p5kVOwTqB
eK4lGTZOuPZzR7ixCNRVWUAlypvc32e9Ojd0aoHtlgVNbpSgZRfzRLsbWry4yPz8IYEu1txz+SCB
bCYbpzZGiAkRRY64+hNOrLVs1n7w8wyR3aA+Jxk+uL3gLuX55rM/L0BOniGe42Dc9gh5pW+ip9o8
r8uXwIIELLhtXvdD8I9eHzEdn5uu8DeALxtC6BUZ5Pwhf4YoWKOaJu9n6bt+dBJsoQp5+ou/Ywyw
hbw52K6zz+O/X83HjzSmPjKFuGWJSIEvdCx1wHLvOOPj+nxyjVOlX4Xqjl5mqHwwYtNe7W5RaCRx
5nA2O34Jl9MRBF8P8IA7tPPnXVGC83NfOgUoBQXgKuY+HzpbTl8IHUgf3iu2Cp7LKMOkYjCwc+KT
kXZWcz6eJSDni2gmsuw/S88Xu5eRHF3N6TpOhnL8W4/WqXtp1+XnZ/uhZQGhRPVV/jGvrjRuAGm8
7hK+9aK8bheirthKvkreXNdmMHZQL9mRNOvklei797SXJbumjkZkPkTVZEzHXCTIDZd8+BlBOhtR
VswIPF/L9g0KB3sLq/n0CtULjXhQgfMzIRVX3cjXgkSIokGHh7NskbhWhxK6dysS06xHYYJioHun
R6/L43G1TpIac/egqMYqFtrR6twbtNAb7B8+FT07NCaZ7P6sZ2Xd0893uCL+qRA1pFuG1IGd+qL7
SCbzwBbgb4/7L52I/jflGhEgLj6hulXwGQY1FCr4MvXeyIK4IDNCur4k6+XroxY/kVQ3c70YaYSl
VqwDx4Qz2pnwGH4aCGOsoJugsdJIkaomacv2PTQHqcCoxYVuV3WR6zXKLJurTQatvK+cBAc/VWHF
wTQa5ZHXuPv5CLlyKlvdZ11nciaNozc3qx2MpNl1snhO2x7vDdsn9JaZNIPqWBwXWTdlR0uBRqlD
d2CdTUncpw/VFIj1XuNhKSc2Mc/Yy8oJJWzUCSezF72zh/JVY6xhf39UrAn4WGnXDEhIm+iaztLJ
2mXF7kMBfh+mFbocshlITyFkqhaHrVeh4nhYh56XowG69cVeConmVZnYb8+mg9Q7gxtMprS3mBGl
5jksAFhcIVVoSGmFZ1Nri7ONTAXAImLRS2lKKf/Agb9168ZunDfbiUE0Pk90tRd9jVVzqNHMTT4L
Fp5sHo0hVGuzkJa7dx+amMeVyz6kgT1l5vrVyWbn8G/z29duRBAgWZLlMyYIEYqaVqATYqL9LQmC
B5wAKrLKZGzWlO5iacmyCZBF4o138uS7nHUv+zsb0S9bP3fTGmGLPoy+UMd+HHGapIPx3junmiAc
UbCt//ERE/7YIy8EbmGKQ6aWYjBQQpZxgyOqymytHouMmN9vXBMTNT5ctSN1zUwifdJfNoNsLXQf
ZmS414hTCsod0Xu2I1o9AEr7z0zWL31BueikDDJDje9/s0vEMREKHZ5uwWa23vBtsZUvyGyzWWto
0Fd5ifRK42QAqtOvj0gK64vzsXIUm0OreZoSyOWt+mMEHZHcRilcEI/IhsuW5yGe8MiDdyYqcBHV
PhoZXqOWyF9/0i9zppUx998Zfebwl+0ors5G686fWDLEobXrsZiWlABmRaGShx5VwMLGp5OvExKG
cl4Iq3MVI10sjBiMLh8q/EwbZxCbZxRHpwsrjY3oh96EM9Fz3byUYv4vYUQqU92j4nV+tmvObmyy
ktUj0Wqqa/rz2drmTUeDnqIfP0AIodYwAa5qoBwGhnTRaqANZ4jmKoaW/FuAxTMu6WNMotlf6l/T
Eoml8tHc3sRHBgz+fHJfb0ZwO/3iiyCYVjf3Csjhxpg2gkSni8SzbcCflJL76oqKR16FxmxH+P0C
cVGT5df2pRdA78H+uZ1l+xGMoYqFBQpt7mkXA2cspZMx/wshVHoK/H6F1eOIvIzUZ3UaXVfv7lAS
GQNLgsocvy7P2athLUc+jD4WjXuiugqBaSSPO/AqScxrmO80S6imDjr/Gutr3q8tU1NoPTt+uuI1
JgJPvfp9X4mjKGsTwKBZDPhbmMkwLntDnm96fNco3SCi7BivG14WoPyHxKlRlsjEfU4OgvkXfQ5J
omrDbt4uVrr9HkhoxW9oq/6mnSKo83YJy/PLOu+c0Xz6crdV5rzrB6KYXQhQI/ykD9X8wolY5jQe
++Sfit510Mg3YTlMGgNV2kr+rukLRlf2TvBjQUJLl0K8R066bZdWViweVftGH1Tcu/dnMSuboH5E
RDX3LTGtVTLMtY/74jspOz95VyTSpOxk5SP1ULXkRKTNlcFaZTx0ROm5glbisgskw4WDxGFWzDlQ
oeVGNQkNnMAG1GNuG1IZ0ILzmO62K8Df9sBbIP0rzqyznJ7x6mgZOD1smcnv4+P/uSr1SVYUUM99
gO5eGbu4A6cBptg4h2X1+9DTxScbhFJLHj2CbOi2/nYq21g5YU5TqS72HA/O1RSBvHBypJPUeTm/
uKxQ3Mc5009tZPI6Co8d+QZNK/cV0TxrRw6s1IwmT42OlkzQPjFF55BstanbXqKfFlojGKuAaNBV
RPw+4urTPuuTbc2B5otWseNNf+K8MOHx0wy4WDBLopQeuwEgtvLXWmhB5r935ZHbcsDT+X36sJ32
nssaGSU84P5s3OOWLSzDI6dOtVfU0iNh5t4L5AQF7ou1lZKo/c/b3yqpFzKCKSyVXWeOjHTpEZtP
PkVS4CEY0VQy+OjV2g5OE7KblR5kociZL9whCRDFKR1WFScIlmL4j+AN5rKWEyJsSDaa4wKkXT9C
6BYcvKaX/Y7AJQRBkB9D+PL6QRqnSdUsm5nLaj57IawYbIeNPr9tNtQgwKlfRi0qodiLxkzOJstn
Q/GrdLBoLbLo2It5Y0vPaP1ogO3lxIdmiF83LXWo8wYtULHUZx8m0xjjicbTtCJO4/+l0EGuG5IT
LTVOrPfKGP616ocewMvCp70ksIFnilJ26zipzRqnSZuPsOrYG0UvskjSCY+sbBAU/QVIBOeN+mXQ
2JZh07LCbKylPy11re7OJcP3y434SlVxWbdf+pLvxV8Z8kJlbwxddMSb7+3RCeIC4UCwkMEmq02P
RVWSQ8UoHo8JSUN/+WlXr1qoiwM1ZMXUuh9tffyFp3l8yw4JxvwXLCWYWop6bdphgGdUBqNWxEd9
8TOO7RM3sC3+DYnTvVdWe5hsu8VlSpu3D5AdqGwVuibPlzBV61+kwDMzdKTwHP4vLfUOhd7YB7h+
t70S2igvuyOu8ttKAh0vbFQutavrCFlKGrqsU1mc42qH4Wrxff9BK8ATHKGUOEWltnhoqxdg8d4o
6n0g4MNLQlXGHWaY6gDVOhnG0LKSZmZXUBG2Y5SxRd9behciw+a6FmZOz5A9t76tgU245G/mxU+v
VDI7hT4gozonjWS+q+DJRt9buUTQvg7QelOoAPfYlJNF2prRuQa34Y3Ho9zZQnbmfm467rLa2ZGw
WCbZFAAcxRl/xP8nYoJPanlqXCClQpxkgUcsOmVfYccYOvQywrT/DeLwrO97SAyoQSK6rWkZVnEB
eTAajZ/SgCR7jTPhUYpq9/zb0UnAdpGldr5yXE4jfvj+aOZc5K+VxKIfe3uW+lrEJuNA7vSYco7g
izuFDaxBNt9JX+NiT7mM4P1MrhGFV2fpcSX265Xwg6nuigOy/qfPxUqykQVRtO+UWq3qR5v+G6nu
0KklfLegMZroTq5Rzw+ZHVb+ML+ZEOLyWu3muEPf/yM12uZggHtXyxjG3/rWypOpW0DVa6mxGGp6
f2e9O6Q4cue3sJ2sIuT7kieIu0djiOi9YBRCoQ4kmaAxVWkLMHSbseWNRh0c7WSW8+2AX+ORk9GU
IaxZxEFzWZhDQQmZjeDRoU4lqK1Ghk7rdGMdByN4idhzN/8PbNcUiXAiigLlxTxBtelGRBSeUJzW
w5N4tXD/kBmSjvPLBspOq91K981tygTSbO5hWaj3Rfnz05H7+YbJ0EsU9Kq1l82c5jmhQDzn0I54
4/3zypiSAn7AxaX2QFHCQ4ciLggh+nFtv+pGtbtMILK/08RbbD8QT9AuIEIE0uiKD/7j7xpfDwDV
2yfls9lNmL0HR5/CdrmJZj4pytTDLj2MYLUgROPID8QFqkKD1TguHpAzMEIqdzZd0eaROWzHX0L5
M1OFybfOxotc+g+1H2122Oo/REPCwbQYikNS05kpOaAsAC3CltdKtTuQY0AIC+ha5SYC0FbMeFZt
6cAiyJKd5y291cRPM32PNMZysaprPSlrq1GK0c32RlrVNEv4O4Z6+k5COKiGmDaBS6TwSLiApMLh
LUOm/vhxniMtIWrj98LwPg+G1vjs5JgcZ1Y4fJYPqFOF5SSydVAumEChLxs+0PNR3Hm3UbGYf1VK
+1iRgpUDuGDJxop1hc79+dTVIUErTCxjbBnm7EnFNXFC57LMWgAwxxg1d4drsSsAv9t9l0FOnIUN
cUwRjt8FK/0kvPtLSo4OguH8ogYphV1omDgm7sQ0mNxsnt2vKXFVjkdcHhwyy7w++kqF+biLqeJj
QO7tVyF+3s9KAn3EpyCns/NEMZktEnueIo3mgUcSMy3Q0+t57bbBzOeiioftKjOXVf/UxbXrLFr8
7OQOHUS+v65TUhkkRJeW9GWusR+Zk8qNEuq8v65itTZHHiDkAv2bLZ/jk2IJfev7AOgo28NhIfCL
hI90O96jOHUxKp9z3XMyeu+vThZa3AheKt2G9gS0G3we5qp57V6xbuHG0XNn8Fu3wla3VzhB+xJM
BmA+zhUZqCLthbMd7iofKs8w9cCC+XzcAHaDy2nWBMfbAYvGIY1mYr+ugAfusFJng2l5sc2Y8hLY
8tt2UcGpUe8XPXpQVAH5SrOubPinABuFu7WmaKaiwsRDT6oF7eblfAcO4ZFq3lpuw1ZnDbyZJrPu
UJNxT1GwS6ITbCgBf4sxWUJhOcfwvM7nvUrY3bd5pv1Y/FS/lLt2on+wE1+zXunb0ftHYmcXS/ZA
3escOrAiRoD7Ds3RCnG2oOlKpsDVZbvq5nyvdiy0UKLWI8tPncLak8Oa64wNbHx9XHJjcOijaVh9
NB+b3wfk3+BwVob0sECuOHdlQewLiM+ELWGTdoR8DPS26qd/zyU7EjU4VT4ZmA7Ezy32EagGSwR8
euAQ1S0ozHrbJkfovno+qEqO6MHu9wvejSN438K8+jRpR3GX5msXv8ZV8Io8uisKbteFCHaUCom5
iD9sRRRHk8sc5IT7MDRP7Q9YACAx32abCgj1S2JEzId47fjDQtSfrQ2K1CwV5Bzi5boKEAdEqJXC
xu3KdUBAXx0kQZC65JXfgoo8hCEanO1enhYJieJTAl2l6j4vVSvBdFocX/7dqbAUEZRzCn65cmEP
3T3dsFvuARw06sJykDRfHZndYmLwPU5GG/5cCRjPUrNXERAyrPX/COHKCrpVVw4G51+5QQUSstV3
uN4RtG8u1lAhnll9A5DfPb4z7LDXUUuOeFCLNKX5LUg1ULKrECa8S7c/bagyXZJkbhJBlhpJ2fWQ
cZkXeeL9gbHrDsQwghIWAuU0hulU2fQWJPG/jYGwwkGU0Is9Cgal2teoL6a0NdmCIe4kK4iRiYN+
Tv/i52qQSf0DHdXDIii4sJJNZnugcYpjTd5wLIVeFx9PclkzAeHeGNY0BjHPaclD6Q6U9eq3tVkQ
yaVVck8FHwuv09Ngyrrdj6op7q+adiddT5sR36/Rybe2vj586+ldzd2W2otRCSCv0HDZEL5ZriE2
csyBs8RA17cn9DJg34dU5lIM3kaU+rHjNBAULFmj4MWN6gf2EYqvSLTbYIli57tvx7ygvcdVcxId
KM8m6m1wV2Oe8+B7RFYLVEDT0heqmzBgm663Tp6/k5IbrqzThuqQZ/Q39NQpUB+t2NgDacGM4cNY
SNvVtZzq4mdniJ8VgTW7eIub7nStXXtv3T6APe4ibvhxpkKnANVnPNp5dLkPjesLOkyHiv2tHerl
ic6cicRVv5MVS8OZUj17N9z10wpU5Em/HoFxaHvz7iImMS16KiinW9Z6aF+t+FMZkclKnBSG3orr
C0WFH1O1Yzi/EepiVhwA233fD9ox4xvF5RU8LvyC+nHduFXngRLMlyqCe1Gx56JEDwuCfWIkFKMI
JAIp9/ksuTu2yw1XBkuISm4dOc0ybYbK9XlHg6py/MiQh2GgQ2VIAp/bgu9ZFRDOmYaBHALYf1em
C0JMDMAil4rAlM2Hd0yBcueBlr5FQWFaXG00SlCIGV34Fq9XMPp9BYizFos/2eDYltXKL/82br5z
79z4cMN6/7yzDVfwA3c7eDUdipP6IWuF9IKfCwPY/U3lMoSwY94g+fDKoBi55i4zT/zAlTWmjter
255UPlR0T51Jl2xqFwgBRsLY06HJ2VfKsorqfSWcbkqDMyTX12fSh7oiB6EFP6HvhnOxYp3ek6nN
v6mxXBAAJua2VwtNMO5DcWGZYk2zvx2ZhU5aHEg4qYSUAf/nAyfDxrAqIQaeMOzH5uXcMIAKvo0H
I0NhazAMtdNn36Dj/tfG8G/K/e4nxjyAWr31wW3GbVBw4gd/Jhi+UfidvhSctND1u6fPMibhoXZ7
o56+EzKrLtypwuPfVu/ktCpvsTRoEwu0UsnX5bdTY74+HcpImG+QMvZUSrXXa6WOfrzJe6gJzzuD
VlXll7l3VdcbJswZsxittb6pOX25VpYwgZLOuD6/hpJguJ+3G1N7eMIFh74iQI6gD46uh/fpGrZf
LbYYwEeJgJxN1aBzUUakIHMaRwFaRXdwKn5WuvE0Lt0ePezApLBdXOmAK2jLqPnMSj6pvv8msLRb
QPGR3B4kfSZ+EGHmlKMkvqH2PW8TtqIwDfUeauvRTpoJWeOnTdRxYWun/wur3uUb3AS3GYkGWIix
tO3oyRPAioVCJl0daH3+DxrWhZGwhdMry2toHHvSIw1Kw37X4x4uHb16+Ejwy5Q5G8hoBcNfKCB2
S4hsCIHlg6z+yQbo8btHpvwyr9VL/+wsGRePvmpQHtUdLs6NZHVRdfQIo50b9upJpdUt/1sRSOJF
JM2Vl/DGLGhgKm2BVOT0SvAOLOYW1DRCjlRYB/YXkV93fpBCBL4mFhy9as0jtWwW4rdtR2KKM72K
8n1H1NahfPv5PMMPIxE2CH3Cm/TzvPE87IQUCEAbPlBvKUJhO+caPqUy70kdt1XJjwtuTsYAeMBP
FC+m9TPF6cFJr/c0yUqqqClQtmdAljZjZQXJ8ly+rRzT9JE+3CDfNYBwJrG9YuL2pnxkwkWbSHvT
Oap7Zy3KbXMlTYlhkThphvPK5Lg/4oeCzEMYNAy+nQ7Nelo+Rqad+wvPd6MvnpnunnBr2hteI14Y
xl80E3EqemlV3xTk/jKrHGorVwSyeZpmyl8xPJDNbSvYcMVeurBFqTJjlQ5RRMDLxB9jdChjawNN
YoIDmAoRc7R0biiTpdQXGraTxJ6d+PX1oGJkQ1wErMhcvxeg/6tCx2Apc5uEa8S2HXBdqopAxcrM
ziuZPOtl+Oq8Bzs/16OkX4NWwavfqa2a8Q2tvyAPeI74eT3xXSesiDmw+MDH7qUXJjZEvdt2kf34
jlENjowQ8OGVhWsQxMwaO0367Jg2msFznT6o3Sryk15j5Dx+qYP3pibObwEfiJOsaggQ3U4wjUmD
KBTeaGmak5Bw13qOkPw1UHN8oYa8kpKYaOTWI1JWqYLj5/9Uy+7AwqDoWea4Uj3i0glqAzE8ifmA
ZbZxUxIDC8RRXugZcL4tK2X3MKx7q3hrzUrXZIwNfLvqTzkCOoEjzNzO1kHoS0dptEFcYWBRjLUe
x6l+zqnq5RLcwF65LQRhSFyHr/9NtFtlR6PlZMQMU1KBB4Bn4mu1+GFaqrCHF5HCyhi/KxN+Lf4I
CVwYc2pGQouR8exOmPcPuUq6yXR+VgCQtB6l7cAa0Qnoqya8bOl4+ThLL2d9FgncaWrmQQ7arGxr
IG1dkARcVXb/DaBDlMQnN8YyijUxmTw1xFbJ3vQsCpybDdQziPivb6gWRJgpK+OwfsDNtj2d7XEE
k62XbKa48o1bqBSsEwyg2Skx8o/QcXzdhf8E93/oshCxF9qChE6D6jEshe819YfoQ+H52yxYAFJv
VnN9LPVk+vwC7iNdmGv94jvazLo6eixQHMrT8cQrVCvk/SrVccDtkT1HC1pOXaiklrLhQzpo1WhP
P0nZ2U/bO3iujAmBofFUc3c0egZYLCUFfUYOVKwHQoa/W/POr13RNIcrIVwFusNdor2vPLeH1L00
+q4jYLbMCZL2A1XCpk7U+oqBZnAAaF7MtyKpRkiNXHWbVsC2myP7dsJHkwG+uOW5e0fBvVy8/p0u
iXJRlJIQaQh2OnCTfijj/lTeOlhlOQOLX/P8zFuGU4BQIRlqECAdXDbGw6Z1PqkAv9fRAfqvgb0A
YdCHHqbj0CgGV0n3vUp+EFmFxsx/0Pe7QPyTokfmLrjAndlrtPyFR9oXhTOf7OLvaOi3xiw8u/Hw
53mC2wnr0AqALWRRlXg67b1d5vN34IT2jNLTbXboCW5kmNa/8RVmQ8G6FMinnrjPAtlQuNoU47n9
bhoOnlPTq7tLGrX56aJmRg3h3u80WSML+3gyK2z4ZnWbAe+dtDs+TUga5cDkAXCq/LRE78ANGdHI
JG0KmhCt0/JXtVKoZPfUFpeN9hcM0VGLms9rNC69BQaO/XGzMVdqFxcjUjhT25ltN3X3hM+bXxy9
ofJP5fnuL0Ax4EOd3LZU3V4Bc++pJmWWOXvnJiowRRNhBys+5kRfXXTVDbknYqBZEOx7mgc7r7sE
ieoyj9+yBlN+/NOtaShFPkllsHmRcXIp4LuNFnieBVrz4DNjRfqi1Z2mDlAetPX3wk6K8WNwpTEY
CSFtNVfas5hZj6gzcI7x8M5pPAHzYF+pHPDZDTV/OnhC9QVhQCRoKVq1LMjKHB+dRZmo8VBzyDon
l3Uzl0mQEBbdxiHmOKLTBjaSRbITtaZLfdvhew6FNVAwSx9kgS2mVDxxTnovx/Ssj91FYoATn0RP
3Lqc5uuPPPf2okKE3mN/uCvePQhR9NqylJXyLGxMw2p6tzATk92nFk4PfT3mo8pHPeKYGphl7Yfk
eCoVMnnBv07EuA3cAg/iqeP0CgN3/Ep+Y8q0ZVumoYIxxJcs7SO3ogxnMaQeGJ9NoaFFKNskO3Qy
e82dG1AVZoUk99TuptlGsLXbsmiP7s1jC/uO0oBi436XPThmPUnBn8Px47FIxvXwu2ykv6ursU0Q
v7nf8vMzUY4DmRj6+Gy8GkwgUNI19wKD7C7H182MZSwqsGPMYs6rpqJFPZebbeQnv/kWCVb5zTaX
4yis2buctvijni0f4gfvMvdRm3HRUhP6ViIifpfLjUqrJnfhqYP56PXuHYzWVIHsNZf3Sye66SHT
8uTecG20urWUTWmfluRiGk7l4GCuz1xIAmHqKZBeXNvXlaUg0P45ufSGsLidXt9rfoYvDyMyLONI
Ms6A3IzXCL4KDg/B6ZXKu2mlht5jXffEe0Al5LXOyu5t7RyJFz1UjcVfyqkPAtxzxTW84qew3Ftc
He2aMxs4JxzxnVyeHkDIS4aqGTe+GxWbeGTJnB1rBgjzh4bhr6ySsE4EvRACY3H1gFCoskf0/yx4
eCpvhrPyTNKFQZNHSGro8IFGPF67+Wl2A4wHAakHMnTKYr+X/wljPaXh9SGBijUv6o7zEFJVZa52
DlL2FuR/y6NePxhnkOH5oOyI+FOundc/7oEkZzn0rt8nsq6BFMxCnbhhASceVWpoZRUKmZJOzi9I
hBSPNWvgElW9zH9KudMqJGhV+ySwg/Dq+HH32AMTOuheVuyNkrK/MKyPbRDIdjVxmCDieT3FWg8H
jGpWCtfgqXUom24TPI8EdJfkt/pSe+sVNDO7/n8jN8Xde1lfYSxxYiNrUMdWhl964+fQZyA8MslS
WUUWhGa9IrDsHcG5TxqLPvkHBlU78Mhxc0ZEzUNMPaKJrb/oBvDn+LwtGrai4yMyBgvGZZauGApg
n1catzuwuysTjf4Su07gJZdNWq9ajzlX7+OIrqSSGotDaidX+qPc2dlb4rA5b1yrQMGWziH3Z0aX
pmaArdFCqxF7V/NWSd/772poKEJ0E3iKFaKWerULGlvWCNXhjfyr5tJAKPbzlonbrx0HkzBPBKYU
5l/RQtV+HeC2nUxY2tNtSbxFfYJr/4dQ+UQzS9konz8DMozk9scwhobJ9onavWToGGp8Wgy0C+Rf
KGp49WkgKYzotVcoQCBCmIX8R2A2OfdqWcwCsyxVOGhzO6goKWo11JtHzd/Ji6rsVIy1ziXeCIkT
ZNNEzYUhNKwMDXqqiStpwG/w+G+oZlG+ZLFV6AbcfH2Kyo2IKsp+SWUx5JIaoS61W7tDcOpg8Uzp
Yavt+j8nTVwPcu5jbeP/29X2VCQ4P4qGrBlQcb3S5QHyoEYGK7Ygzqya0C5F48r5my4DZ/gAY5hu
UNo9NYOYmKvgiROjCAY2gjSa8p/qhmaM2NO78MVLJH7EIUe8p/SVRvIyYfwuTO+arq5gWHGKLHcg
xEFgZPjJ9Vw/VNniQ64KuYTCBFt1/kBqBdapzMNiZHdTo703U/F7BDQEnOKP5LPLMQRxVzZTgJ5d
HDIRFSidyVyBIiQRM+o0WktiRK5ZBCy8PugU9pVjHulcE6WrJDtiyAeVY5PvkO/kwskUa8BrFu3h
SeLDxCEXt/77JOCjVWkY8WoCE/B7skflXCzt9aO7Smady2Iqr3J+OvBN+dyU1pO6rzr28FaLKhMo
FTQgrcZuWtOz5hckoOjXg3RuZ/iCIUaDYAwlyk9NdSh3CO/3IKTtQ9dkdd+9tGLiOA9H1Z7C4jZQ
yWsrYNoZpgurLH6Su6y5mCrSu/tia03DzO7hr8iaEP/YufvPzWf6Fu7yAPXPa16PiaGCgI++K7u9
S0eqQOscI0Y3bedXhLnok0dQes+gmUwccvrZVN6nQvpe+nvA+t0E5TdsO6KTMVP5i8goa2T+cqqS
b9NiA2mKTbX0qouU965lbLMa1z8kJEJ9ELyJLOvWboxZ+SBkQwl/6Qt35ATNalVSp0HblDNSBbKd
wtj8JN7SDl6TlIPI8T51UvK25/7003jw4ixbLmUf3QsGJTrncDjhocJB/KdrUTer0jiVzHUkLdHh
AkZDjFEotTC63dTf19UZxqdPl0xmtNuklKA8aVjUMyCL5uWhwRlNNZY1oiC6xYWXzXgZJYgP4Aju
wMxBOECZopoc65xxuSROG+aUnyO7W7pD+ga83GHGkAmfjXqx8EtTWbKZkmpfl0ZbcC7QDN3xuCLz
lFwZf/bJ7R+wnxWqRbrKqVi4Vh8PiPXQIVHsdobVov8TK+qtTnt2freL8wiItj/7U31512bRwSS/
pWIHVeXmIyOdvIc6oCjrpsnSqHURkpGKnnAjIWTYRtlEQ3KFTuBKf96jheGFABXF8uSwqejzJj+G
jlgCwOm0LIbky4idT4NlJ0ksAaBfIac+UG3PO/+wTJGHZ14vTMrWQXzW2gPHyzb25oNd0cu5utbO
0bWoZRkYSShlDj/2nLCT7E1vh1MFl6N/QWeFLHIr2Yt3HA/Upk6TsevZU3xMQFjs2qyaG3CeTqet
0hN2pY0lhvyOjXKau6mOX30vxs5vGTpWZWXWovdh7ThqB+kL2/7k110HuweLAElxoVRWtZOBui8Z
O3mDifgvF+kTB+PQL55Cyx64sQEZlDfA2stigGmxo/2U+2Ks5mo3xC/rQrT4qLoqcXrzSwkZ5EyH
PdUkINjZzrrgRANi+yV/M4mUUucSiDHHJPLgjzswiDXHdELU0z2GJDIA5Mns91IfN7ur+OhKKjk1
ow+53wrlVRZr2lwN4Yd4VCbzdNCSt78SgbV+01rJ8uuHacC85omY75dk6onCEXdGeVNfNh+NH5H6
0aIwZzWgVzdDkGm57krDsT3vaeLSkMeOwAR4E+gO/CNwvntyk/JwF725bUW3EMlUGq2W2dSQCJrv
xiYaX9gRJ5V0aI9moD8LGuEBIRK1gpqOiKcyHbqpyBWSpD44kXcEXEliWEbsAO1D7SDtxTvPrs+z
GlD1uJl5GNUpvAAO296JwRfKVH7Nrejg6IDeWGM1FrBT7iFrMJIWLRY+nvNf99VoJOVukMsiyGSq
U8AOvLyrzSnkc8Br3D8EcHGfnGNX78yJWQKnS5NvCusnVIR0CcAFP9AqXKiSZ6vw2QCg/7qP7t6r
9DJ0ZgdQW/pZOzjCw/YwZngVJZbdlDC8dHBBQ6Aa895pMYHu8IEOaZL4W/TfWmGThTWwpU0OwKG+
WZ2cWBXM6TIP3EGJbQTtLz8ehoRcdqw0BRW0g0cupu5C74IcSaVet4xot9Hbxo8JMVqPD6h3HKiQ
gDemLDZvVfON2c5aANW4gSYk/1FcLQqY7Czv5nfFmv3wajpoSvFV5TdhR343DHdSkJrsKoWSTjBx
H9T4Ykd00z8zrcJq+bIukpuEUx6RkEVQQGcEUhSENlx52afiWJ1vEAa5T2fMm1RdpLQjUsKELiH1
Qj/lGqNvg2fy4P8zwV2GfoLds7mQtC+vRwKlmMhOrhaiSjZnd1IHqR+TrPa5ei8mDxlmEEVK+o9w
X0LGY++wkNSHKQ8INRItynR1bOAK8KbX3R8u/LmYkwpZJ//EhLV+XJyz8s8msww2+W8BekmylnSV
vjcA4F4I7IdUwKibtjOqoLCvwyHE9RJjxgsXfKQhw4RVxPYNxbY05H2OumwEP0le1l0/2G+AFmXT
8El3vRy9CtwhgoL9ijjgnTi6uqZHhhq7zysoICTQ8xxzjZdhL9PbJPDvK+7qVt/nvgNn8dXt2Qcp
29g/ACRNyd/tBr3ZrFT0TiNRFLzgI2t4YvJoqCReAMvlO2f1eoxxhKRyA6l0nHwuW3hNZQfDy7yk
V+Z4o3HQTZx6Z3ZNJqEIxPl/zrB41xpKor+XI/8Tv3xitzuGdPj8SuZkf41Je+fRACBOfSXDWIiF
BX9v/ggxQNX29XJhaRBTCWdbNGagc55De4cYLC5xNZaFv1Nywt1E/lwUQgti2tBtbOYl64lUNkpA
9PwqPxfurmYDUeTF4AOj/axCNmbDulx49Xh9xS+U+QhGCQ0f7ae3OlkIaChYuZaieKb5UqMLWEtU
0ff8G+0pv5Y8Ej9aXHGgGegzuc3K4Jqa3Pyw08r76M3ts9EaNYHj6wp3fJpV68wio/7uPD6XJ15g
4N2ujte2+ziv2BDU+j7XsoQd1s71n6P1sTWwHab14ea6tZX5OxFC7xZ8oDrdlUMh/eyr7duyUFi0
iS1VG6iUMpFY4D96QeP9FerDBFarysAnncGkmeieNsUQYNjCnl86Usjf1/G4MB6HF98+DLssIRIs
CTsHOS0/VKw3nkLW6460jamzF0fUoHDcdY7k7/yieW1DIwKa117ohbIGFtDBiQqAogwDMTgrIbjB
KLm6WNGKV3SQhLD6BxyShuY+NcCMf5eLr0JET6Py0zyDFits4EHz/XVH9Xm0kh30LjrKpKE0nPQA
6A/WuoGmgu3Ztc/UUelvsTKIjKVMy8SFktSuHUur2StJysrkKyQTGZGf8xMOZ5cBA1RFZOTauC/e
gp/c/FWCzsUVr26DKRlTNwenkxdgGWtFy0xxvpU9i3/l7RQYRq25GWUO+ugonO3p0Ou52AU6XaOb
2FdtMxMoLEgbYnbkX2YgDI5ajmAein4Xt2cCaATsPP2NQh9P6mdVUR5y/nz9+gR6HaNkpcGVKTQf
CKauZRvAVGqtfijvxe3/0iQtVJkq8twzUdagCf8xNLSsYdjz2pG2kxcTkko/9inH/ojep73fpuwZ
sPIQWreAA8wN1NE5j9qzV7x+eujLu6Rwl3UxypJ8MXcLfTVnRDIX5WDoiIRh3ERbZ3B18y6PiPEs
TKBEFvIxkq3t580F6neG/7SwF4ZGnSy7RcVld8VPOCXIgw5mK6t6XAK+vKWmvtHplRCXRGClQK6Q
MHJ1JHfkQoFBTimzEpmJcu5lCaBEt+qRVYv9Z+Rk39lg0+XPkNMwrvLG9CZUZFEN8X/m5EEhCOA3
G7Vr4pxztfCsVfKl6gkqXbIBDwo92omDiJy8hD1wEp9kTTV5JNvrX4p7aTRxePEX5+3VEA+deLjK
nIAifMw2Dr9stn+JOnOgzbr0KPynrmdZasAt2/1jHYSGyRsdE/Ubz35V0+61t2iwL7JIobXMnAU1
fXxkw9VodPPiqyxHJiBag0gNAfbzoCFeffXdjGq8BMoukUVfjMA1lohpUWqL1Z6T5bTghJW3t/Bt
MOVT9oGc02rWzK+tl81TjuZTdOXCrd7zthF4/+RAtvf4+5P3ybMl/xicSTwlvrDBTJzwhrI14jSX
EEufmmVe2dOh/19/XNcXttAFB8s4epjaY+DDzWbu3szZfi7llY8FavmwwbNbOQlu4/uBzQo4SVGB
g7FqdvmolF7mVuQmoJ5UspQfkSWGRYmwUB0Bs4aWM5mICKnzGLfGgjqcmK1saxcqr4U46Vw+Dnp2
Wq+YdW3Q82ANvCQx4sY3yJUT071sVzaMih7EZJGpO3Ky/Lf6/J7mesGl8sFeo2EXnyaer80jI3jk
KTOcS5qyfvv4m6p120OV4FYZWUT5vL2KvRamGDhCAMXaQMSsUm3ZyZmu9L9C/Xw3TjpBJ4ugy2ym
8q3UgZ8LZIs8dRIyaAPk1HS3/G+fzpgLczf+YL5s2Am4pu7rlKmMtyX17m+Hc9GpqD8wdDbPOmx+
AjC8Sazd7IVd+JqM9rJoQT8HogUdqvvybFAxSioGn0yNOhD/E7fpzMrGhZhYe28ZjJWcywbE+5nv
+aspAD6bEJgzajs7DS2DRq2LdIbHUMsoUt2kXlFUI1TXheBaTyDlbCevyGDHNnqzco3EtVSMWbwl
97GXdgSGu47bRFYNEhI2nA8UF2wEaYIonfN/Eivx0GMypBUaCAyuCQ6Y5Aks2EzNvIVU1LAXVQZx
bEpsBjixMz8z2H0zyNIolVQr4rKA6ku7onw6aEBtBC84gJeeFd8I+40zXpERZZh2LiUiblfn4P6o
Iaan8EjL1b2HkrNXTA1rE3ipC3oCIHZjb8iO8DtyAiMUKLn/zQX/Rrsy5i0uE9yjNmBWjGYk+6YE
1P4CIY2JnDjm+5nFfXtPzFJzWirEF78zZRrmtjxKPis2ijA1g3GKnhIqjxSrJ5TcreKtdCmVQLkf
wy/fig/rvcfpegKpUcpTJXruCrLTYv27T2vWM+m4HkeRIw4XUQkKhCqhJ8DFeXFcP4782w6NLqeC
YtiWk7RDOgNSstH4FjGVOt3Ks+3rY68MdFzOJV9JeojM03cK1hBObFkIKlfYm21aEPni1nJMy1MO
a8wwnVH3ApGU2gxAX0nAoPpcTOwVX1XfKYpQNGXJArpdhbHYsgla/A7kFy/HOTR4mTYmOf3PaHX8
yLrqKcnp/9oXBqaNZYQg4F/0fOYq5cEKLZJSja461TNo3POWjxkjX/MG3DwZe/iQM87mz94SPbvA
PG2rRToZOvTnd9Cb5QYwvxO0FYkx3EqTLsWCM8zDu2tKP/recCMKSjn3EvHRkwiKsPJhgD1dvIPx
X/oMMr27vzrqCPar5Du8BKeO4B7hPazKq76DW2WadG+xkfmsyymbtqX25g50d3+y9XEr0tCFvC/8
ZaeLQL+oSorBt6vAC1AnFQzYxnvj2nM0viX9/7XwpA9PeA6R8lPhDNhy0G4ARboesWvcqt1qOk+S
PW7Xynh/3j3yGBw2Ua9sG3OhEN5h6jtX6DjcVTh10bZhIjma5wDDOmlijRAbxuMOFdD7i/tdXGrV
U2GcBRXTWnRP7J8uOzW0ELA19sfdsX699+cUUATGyY4xpu//KVAdfAmK4uxFb5LaHfNeZ0DcO/dY
BM4Ga6XrnY4Gk0QnhKAk1uYbpOUdOKCIC8tbYgljf72l+MLtw+EEQW8V/kyM8XMhY0TelU5w499F
SNEhUZ6VGVtD7rvgQDJ2pVjYH9LHAR91s8o9gpswW5rbSw6LtF2dZmaZQkbNguOFzwVWQSYC/3gu
ylIAtjp2l54htPjKWa49MoJVadH3wp8hAbcjD4xdPRBqJNBfYCzrkPYVWBhdrYpykQoTi56Snh8C
ePtZknslm7gBLVKz0Bt6yY+GO1q50ikjWJg3JFKzJWnwx8I5x3qXyNL6xSiKZIJv/RDdIihdTtFo
EsaMiMSyUsiRreSLxQGK0/AN0bZd0BH26f1bn3jq0Nh71la3X3Hvp61ofDurtpPrGwiubs14/Cib
QF+yrO4uhPOgD0N6siwule/YWzSQ/O4Lgq2aX3YY7DAU08CxSogXlAb1faLhqO1zkIzWnfMbKxEy
jxHn0r1/jYUOkoiFk0EkDqfeIL+M8QfZrmnF0zjMTa7x21/LuCJIMBGfRVS+H5f7RGUh71mxnQPW
Zpdpyd2dFP7j00L9FgQK7YkFxeL7vawFTIhMUo54AUy7VWLIzNIsF6J+/Rywdz6CTSFiQxOsak5H
aHvMaYSyaEinAIpOZE2cmO2v/0y4TaZWzBT/Us00fsrsu8eqmm+IGxOMHZLq2BT3cw8RO7QcwQq9
iT0mpu10Uyy4nlElQSxBTy8fkWNpa4Jk1PAG1gsFw6fb99lI1l9rIKaL3XRoGkZ8EkI0ISK0T3lk
l539oKZRkDqSAY8DSeocfpFldonuQgydQ5oPt08UPv8hfbSSU+IQ8o+jbCpXneriWjRqrris/hly
d+l8bUe2lpkHlZc4JjwAnk+MEdEHF4vVCy9yHIgEA3vzC68fwX0h2+QGmZQVKqIafhKn/7ND2af+
MCwBkZAlWxYZvRPPP2Cb/HkUPHvAsHx527N5VBN/L21GPueAqXgKp8vIvfl3avd3LN1jEbdPr7h0
v+SvYTscSCyJ9lsvcbn2JRRN71h1h/hj+slupEPYpdJ6OzOR9oDK7mR1enN1emlvjkZbpFoTBerk
k/r2aAJBKZsgFZIWEZu0k+1CL3svDdMyzJUvVhZlnaJqX6z2BR7tdgNa0z7fdkInMbZTAjqMTjCw
nqZIHzud/PtJOt/8nU0Na/u3darmMDE79HgQqU0zm3mhaAnXjLylJxMfCBwIKnVWr/I+7IoDdhAM
4d5DkN4Q8y8QQ8dSuU02CVKgX/+cNeWDH/xc2PoW92msYojI12iuFhw7OZoAxrwHKMYy9GVpaOcr
4iOJ4HfaJ9tt6R+Q2dLEwIpbsrszp1AkSihkFVRDQMEe1xJFaRtdklvCPEyVUUCHm2xZMwYB4myG
Zke2qbTJFYi2Uh0hnZpkciKkn/Yy3KOYCX3tf9DD3RelNEx34zOmNOyCqZmPvYqIJJ01kbnL6xVw
9NK9zJ5H8bmaMDBT9+7jPS+RkxsDwrP1xX+UMwfKCd1mnRc9bSiLclT+ai/tjxuvjhQSOA2oPU0B
LxTsV2KQBCvspBE8QIMtwDoGTHNQys6zmYIliDH0/B5iuYitLueViwPeXk2msvoQsbqhzabOJyHN
0dfx09SyWEFTI0V/EBwaz0wM/b2gb2w3DaCKZEMgZjp75j71u3sIveu7YXpWZu1InuPgEkfna6+G
ix8hXU0rG5YL3r8tENqNtJ3UL+uGgY/W3Xj5IJ7V1bDHVZ1LUvx0es2ATNvmXrUkks52LVkZ8e5W
hz1t2yowIX7VwnoDn6OMdywGORNeP/kpCV3qUygcZ80jPnRrs6cKjyfRX9herwE0nv6myyVFs7Rz
+rYaW3L5Viebsdh9+17n3e8Oztt4z/OPgfzED7DUy//UK6i7yDc+xJbfqRah9RCPqa3D0FsROb4q
6qE2Xu04FxMMTWrEaDE/1yKMLohrtyrq5MNNI1ywLfxjSQrfSApUPPBDlyBqiOllD1gnBe+7n2mx
e/ppARvWbTITj+0NtqG02Mqju1pgB7leSyyj6WngvmlWGKhS36A0OhLgk4UHY0ZnGjb1Ajtswsfg
KCm5yVX8gb9D0tj6RoqFn4ZxyTcykQSa23cBC23wK65q/xar/v2ZxbKctIZDs1IUMBdlqmyH30nV
7FFzSGW9W2OhjYgliR2hk1MMRSWrx/mkozd9Otl1Z/SSOGUnf71L3RLmDoRzvpqxtcWgWLjMmFBp
l5uifXsiFnlLL2YrKZZ+3IMNmWKLAcx7OAE33tkG7OGfltEN4ecsai9NmBdwufp8vhwuCCFDA0aD
r5OWkcxNYuuTB7BE05Hs+JilSJN6W0Kp9g2eHu11aeHIqcMmH/DgSQ8kUmbfd3SsJPCoDBY57MBg
AzmQyW5y0R+Rwm1Sa3FbrXgzL0Z/0D35j9276zIKIFrs/+rKCUGwEED1HwY0pUn2PdrU+kLYdqVM
BRJtcmLtTw/bMfIVA5EOyGNxbLWCc0xSWc7Vxe02rb+kvtDCZE8LfnxRz3drn1OwfZ6mkj0Pxo7b
BLy3Jojenkx2q64IUP1sPZTFHJTf3s38oenELLmcIFepB7SBJaI0YCo26I7kFplBKpMBKTfbFMTD
cQq9WHmI6+cecIDQr/CtmIzzXWuG/BJkNeqHtqHwML8vfi5uAwWaeSVi00joZkS5bqYeFKnv1nUs
kLrAR0/iXivb3wRkQGPfOp9E69wIoOXFQIFei09qZ3Ip+6MUII6hJDQC1W3g0UGRD2THlAdPo2wt
souMhRG0rVkXa+liQQmdUNDmYsZfr+oCXuJtQiXOyVzuj3waPeHBI8VIRbF6JSitOC+X3cjEMMQJ
6NehJ2ccVSOg/lxSPAGcnuVuLBvyjl9vRXDm25FgX2jTqXcgFkdTnf+mELhPo0HUtgajeU0D1Hng
eM5H3Hd6UJH/0k6YFur6wE/bBY3rkhd6qBywZqkZLb+YIua/DBbm23Q1T5DkrDhoixl/amsrYnMH
t+2VsDvhiv4ze2RTGrk6hj/OKHkWSbSNgWniw0n4hzREjAQgo4d/85UTQHLvhf/xw/zIE2QT6CQD
xHUUasG26LfSECGNCGdnOgX5uJX5IWl+DcVu+1AIyLbWFnDd4+2ZcqYlFX6ZaYvIJ4LnonLhSMkC
tlAYMR4XxjhN/FTU5kyymQuqIysmnPFtH13mnPeDaMqcynny/GJVfmdviuJiuHJEtRNZMFhLoiXd
daVBj120mo+47EQVvyta7wQ/T8VnCMIEU7DRCYdmtDXrKkNeRTAJ8OqhycdDwmSiPvEBpOk5Vry6
5GSBOQvl5HtuVaoivPt0tnmfMNirxozY8T6F3iRzUaypNiwpPH06kutzmySDXXF+7qYyFA+JmS15
EeKLqCnStjWqXnS1GsvoHB481q76h2y962ple5CQwmzXCO73UgRlzcsY7mmUIzoykiWicTbo/72w
0AN3f1gizAZpuhG4jaH5F9qZvJ227LPkivjbHsbwWV/Wrky0SoKcixXbunsJfHtd0Y6InRBDy8vn
WVcIA3N12bihZHev0u9gM2pqaJduxZw+LJtlZ0PZecArqJh+M0ZtnI64wQRWhtYw3ZJ9BFYaUJvZ
lzETJjcwSGDXJNW3cSI/Ef8LgU0XfhO+RORO/fSn0sdI5rnjSvR2jHho6RGOcEjmu0bOIP30yXAb
DZXSwi8bYbnHz/fU1KcLS9tDv4CGZUKCp/9udx+RNgUm1i8DfBIgjUSdOR90QLkv4FvZS9mLJFan
scP5QJxj0ekxg6H+64Ae0Y0Z2Wxq7rAUc0LGqnHolKE42x0dbEwwGjM43oGbdiuNMqrGCi9RQIgP
nPjVLSJZ4rL3tbavihC3HcfbLNB0VwWEfVIo+80U1QsqNkXvII5jmw3WYLSvCEf48L6406eyfi/z
ID20GHyp7o9slS+MakeNgXjGyJTpZN1iRg3gLtfZyy0OiaXAGolJY/uFxcGPfjqTItDsiSIuo25d
Qmh+2CRaIkjEHFZfo3Wuxg5jTByivfCCUVeFI5E7LGxv22aq8yegzaRPe03puA7t3ZZ5Se76IER3
KUrWLH+RQzMWhSDxva5tiFb3p018wG+fLRrhkHOOxYsUDVJzJyCIkz6Sc96Cn7rn96NCb38lg1zU
S3QyoH4aFx8aeraa0yHK5j6VRG1+MUYrrjyTWn8YUDW9793AdpnkcmPKKyMZ8/e40RnV8lzNoP7G
8xFSkz7rHJP88+g7Cxh3hrgktmWIvfEyg0E4PKZtWqFlTLgQQWlbJaL9GLr6kvx2JW2N+ut2kLb/
IdQr1W2AaBxS8MA1rQpxYT5W2Y/8mv5u8pqt4EdbsHeaH0v3k+5kQy7AE5Q8bVYrhoK8uAhVOUiX
YdMKPilbdmXIWe7RhfkApKWaD6X9e3HXUjOCRip+exQKnLOe3SIVb66lSLl1buDKDJ6Crvdt4KVK
e7jrVQEtJfNkLyauAC3AD0aWQ5PCjkCJ2ughYh1wxNjhqLjKO+FlnLljvLvbu8eySBEUnMkPt65F
3F2PqeXrGI47Ago+O6/kAsJq98boqL9Dlj6vJr2AsYrMPDGWRygJDKOije3H5ehurJ4DpY6k/rYb
jB5yZb8XAI2DI0B7OnJcONdlwMeVDrlv1aEB31ymROWj1JqMkA6YQHTGUFjPISuPWSLwiqoB2SzS
mPELGgOZtyUgLyrKbKbcB2G5d0lYIMLt7xMXtdHqEt8o3M26FEAPkhRFJlsdM6Ip6RKa3cezIOFN
9Q3SvoXt7gAFYhiAKjSEkUZLbVDr2brMKTQWPa9QkBZ7bcLZkoP53TfWCUYEBtH8ZJ2elLa52h7H
+MNWle2iEhxWTwkwe9xYz5eDPHHEbgego4gQlngFJC5uCeO3nvjS38LTu1j7/HXTQV3xpeJryQe+
+Lwd8kcOwvg1xQFRPdaA5Jp7DYjcwVj3dUmhdMhRtTC3EUEZoWx9BzEtEpUSpEjilNpDWQrAXX3a
y4GjEFVK+HHh/ImMm4yChAo//e00AWvgFs9viwch7AWpqbPtIJ85B2NpVvjNDauhim2vkxeqZXHb
9aAiEeFYFabW+ONZ4EeA9wiFLpV86+anOxK0t1DhirQcET1UsDmDs//RoOVSaTD5zf/AGwldaT6c
GsgmHDS4FxBDKLpyudIo0Jud/qfj8LN/8eAa6k/Etg7eQuNZCGf60ouLKPSV/aWfXjS8heZZDJj0
fOynHeA2QYZJU59ILMVTwj66PZS7qQNZizvCf8dVmQGBWnn4qExjRjvtnz4vpRFFZtfGQoyESc/o
TZY/5D7UduFpDkYJkEaA2CINMRWU8/Wz2iMjqa1WmB816KJ/iNMRsXVgdAZfkS7VjbVLqGKLrc5k
0kThA2dfLN8GmXj3MRG68bAF92CE0+FCQV4cT0aAozBV/lHUwuodRYK+ie/O+35PNf/wSu4K7dV9
z3sOeIjsxYYvd20U0GTFt5Q4MddFxjmUZhgeAjHekqImQy1yXyMWQZMaKX49IPTUVL/Rvn9Fk3KI
Zio0qUUrlU5IzmicBjgBdGiOT3fWVXywzOPPOe8+FvqkfQmitRzmSn3QZT8qaYxX06J8SrunhTrK
v4BEUl0kbQWuOIWNZDm2iCP5HKOhHXp+T1IZ6/80QlNgXptCR6ZkUQwBTDW/zk8q3bCtAKSlalih
F5M3JnlkynXZ33HOrXuFWz1/BZ3aHfZr9351GW5MjFg1T6jqA3j4U0VeU+08KYB0goHJnB3ab2Vl
8af7D+kIPQDQ8AFse/oS1sdXWy7CsmtI4Cuq67R7j8isscAmRcvZxtjG94wi5ey6DsvKZQL6AWzx
yJXpW+WmXw+FPlktPC136H6aefNytJv8eTdSNvYpWMl4Zrw2X6hLGGmQVd7B60ZVcCNJ2GcFp8OJ
6MvSGRP0muZ92XUPvZBs1X398EOls8e5CCT0Q4r1vnZ6tLTTxcZlHB17+WAZgO/FLk+xIXYKZEdj
1TT+0L1iqvk/2rervMH3yUGf6XVQZFavy4HNECqaW9QHgsGnQFO8IOi55acUJRzYGYEYCoVJnvNf
QWLIcvoh3me5uIVIyfsfhNLU2hTDZExd9/sMOVHVHwzerdZffeqfAOKnTV+V9aomy/8c5DhGpT8i
sbA1WuuhQlD7uEivjnV2+M/6ZABmxTf0XVV8I8GU61TKvxmCCF9mqypV+V6XrNmzuAErb6xdxe7X
NekMmZH+GvzAuvm0fhs6dbif3Y+In64OlFiQrxnR2lzAV4UJwZEZeB4oUUsN1v7gv2cj4tgrDXx+
BwJDjRjyRMcXbL6pF/ukNOENAERTg2lXx4qWyMqDYGmUUCbTtktxXR5VgwWAVaU4WQ5hA2N0ZZY/
bk1cRVtA0d1VnvvdBj1wnuLQZ3lxxbbfdf6QzMiWhT02xVvwT2ZzkOxjLpd4yVmCl7Pl6MRKxjrO
CfHkXL/TEpzSSu1EGIe0LEzS5KikaSt/KNfRgIHtWTWPOqgDjhUFA4WfKSrvB5uAzv9BehLQvx6/
3lzwVT68NRIsZjeJVApoAq+IpnuMGU1TxyDYLRLJImqyP5yHs6wQLxBtisJEJ9IEALOvdGDOkLuH
MRFe63bgZEjm4Owr4VOxdaAJC9dt05O5G46LbngpKFAT7OvMbEJgl3UgSrsa9xUipPHQvOnfH0yL
D+AxqE4mUNE9FqNE9XJltM2A5KGV6wVa/mBCqglz9siNBjlTOIPJHLuKlNdoRYCIUGqhc3Iawb+y
ZYDBe+dceZobINdYZh2DPm1BAd2U63qHrpP09ebrHr7p1GR44SHdWn6DCc0eycHOLEOwbQfcleh7
BmpA2LQKenTUYFNr5WEg93NDVwm0PI1vRz4qrvEfqJJcl92yKTEKcuEwHTSlshwLjpbTYgzz6AR0
INatHiYRCDTzifgbEACeN/pfYJwt6ii2PMzd65RuD1ih7YqZK9ivT1aeb77BurpT0hMRp3ZNBUmz
iu77ih6B65xpieqU7VJQFQgfg8OoyyCDL/1pxvDEbhCrjf2ab5uney94pKr7cxIz/ylHq1StyOk6
hkJmRoG5MSydf1kRcXVWghi5aJIjlp18PArITRvh0wMXsUSGYJbfP8GuNJVWr/CPzLF0kV86tMtn
HKnetq/JBadZ2kmjSbtQ4NhsUZTds/N28DpbV8pUmktrM2uKughAPs7fQQoYA7nGhLHTBxA8YjII
aEfU8i8B8940ybUGdmOlP/9fxaPrYA99x2+tCubG05e0DI+TdKM5OC1xPvbOzJ2YzW3yU5jDvIWt
zgmEOXtr5h65iBFCR5Q0NLQkm/wieb02ihlKmHFar3rwLvn5ksDhfvwJRrDRsqI35ZDAPIXff78+
Ya6N1L+lOv/55az0zs8yAje1cTarwHNbv/qYpeeI6jaAvvgVpi7t0uDaXt86x/RGTXc5VjoYYhkv
f+O58wAdkk+KQDBMzPZO2dugMZVVSEo1wmlWV1iQow/tr3Gr2FewTnLK/NRYv3Sde9XXm7rqmMHg
RyWCxRsz6HcUSHjEW38/Ns01Xg6zPRO73uHJrGIQdKPYFQa/MVYteF1XZgFtWZu00aPN16p8ldQm
aTm1qgx4s40FwONK/orlnEJhbuTC8Y6JGiTeBp6mHIaDp4KX9pdO1XThURinNgNmECV5Ng8JWtdH
DOgGNGkoUI26wffL4uDUzB4f3HJotAiE+lBDg2qjPuQoDQ+tEWt5fbZi2amOF4Z6bolWHjVwernP
wS8k6mfHeJkcaeYtLA2/0EgYD17Mp1mkr2kWK9nB+SDHoP64nF4Sf6l7wzH/J2Bdp4e45zfmDSd7
IYdPFyIg1vG/UgQr5hDjrHl7nwKBAX20rVkwaA/AUwpMf0aGJZYpBP5vZmnBVXXfAipzotznr0nH
Chjht6SU1MHNBXviK0tv94zKNXLnqE+KcKE7A4bHJks3hdzX1vjqCZy4UvnSR+cd3Fo0Kk18pv8Z
wXN0s5sEdUnY5L+F2SJWiqTHXKWsOaleQdtGOBdCXUCudJzOe28WVRNS22Cg/MGrsPKj29H40Uzj
XWRhqV+48FpvFFlBg7V8yyevp9SQv4ZMJryRQKVjd9pTsNT2UxbvA0Za51ZFDV72zRPC45t65RuZ
dmSDR26fGXqgzzkZrvuLDpVDPLNeTFp8bbLGSWxKQCMjFT6quLYWP7JqZ2bZseWMGkZs5SbN2VIC
n73aq6HuEJwZivNAF0nMOJ0bkudCXFFLyDOACjC8C/vyhcZ2Oi+oma75yMsz9MpMyt1YT59+Tlav
cyuNfBIv8YkIOBce+8GBvDYDE6iq/g9qBJzHnFVLpyAmmLrow60N7ivlbc1PlgbSdmSKzOwIkKp+
xmxJ25drhzDdEqE4CuZ38gx0vmvzijtB+iFE6wiV1/55qs595XVj0Z38YREgab4oUVJIRtW5y0Rj
pqRu3TMeeY2SyY+lO7DNFwOhXtbrEGaOvZ1pMnVUJYNAVYczN6PFM4ggn8lzbNicADCaR1a5d/ux
LEsLAw5rU9/bS9N7ObHw8dzByC9883qmhKR8nLtGFoAvbhBvJhbjVETtzVUxp1qoq1FSmxHl1Fdb
3or1tAp6ViE3b4jOznnSgk6NExXVIJH36mCGyLSWumom6VfdJPcedf+bFRf+VB2ilB1L8T/5ZkzX
ud/HhShdWCkeI1HOGugxy5odMxtLq1y7mGTj4QeQII73YO4/oGR8/KTTkTr1OS/pLsyN/mYgiJya
ohgT/KNBHRo97TNEnJ/HsDVnAgXVBuyJLGn1dAOIDMiuvY/iOTHER+QZ7EujekApiIE27GHg4bnF
SPkDtVpDbVwgZQ3oAeHw3xcRnaGi5yUKaExT8u8IeJ94XUH0oRfz9QDbpIo0MICdSqD2Y+gUBGjD
kDpxBEoiX3xOaLEsm8GbpQQbsCg0IyGBTyjMmJo7jYir9ZhXLARfvDO8qeU9DTGzZTKWzbUSD4XQ
LXjYaaaJjdHZG+Wr1CGMw1K/TNG3StpkIe4pCjz3Oi9gbZ2lGYkpbXaaLHAjool+cP3NClCHjO9f
SyLU1+0Ih74sVnrhqW7gxzaVVHn9YA8xAKwdGnLuG3qnRqNYiYlCgx2Y1SlH/gnv79ZE0pnyo3iU
Z+NPVIf2IRjIiQeVcPZGTXLTYUROevR6nW75xXJKYtfNKK3RvPtDEDAgk4LRGr3Tc844Ofrz3VBe
6wsbr0jR1WdK3/K6QLS7jhLZjsGEcaFIn9RxG5QSFuDRVnMm7/9zWFcAqVHTUJT8145SHlfuFcV2
INrtMwFaZsBDn9TCMLykeMfOUA1ujs2pTRiSZ2+liHOiRBLpsUrzrmOoXpRk28ijoNWAbRTqgTtH
DMNP067j0T0L/tQhRd1ptkv74F++usdReQ46Srv7oEfHNOnUG2+HltDD71ZGSiq5ie+8zWEySq9o
fvIxbjTmetuwuU3xLp+3+77tvLf5AicE2Iu9gvQdQyEQfxL7mIKXkk8qoqOf4Q+VKQ9OJfdU+6M5
JC8R/HAv+w8pPJTYsfLZqB47q7ERfULOLoqKEZAUSYd5KxHGSi39j/i6v53NdDqw2UNiIKl7oPPl
LY7OBFXR5b4yE6vmhk25Ejm1DcdAjvfui6nWcrzYW3cisJQWJ1rSFo/D2EwHHhJcLVhQUIVi4nBE
XqmFmwSHmNIxlxcjH63VICw/Ajhe7j+Au9ZY5jCOQHRXQoqIlx0nZbr0P+l+DpR6twRY7Yp9sDXf
OqS6FgB/R88Sq7wSREPr8BqNPBlyxh/KMDjOQRtjL0R/K8B9GGAYcTUkc9fiMQTPFH5FzoEUrnsI
F5/Tqbhn4b4ok1tQQ2xNlQ/zk431Z8fIWuYxLS5qMVLlGzVRysM7BeJFUzlzNvdF5oUywB7Uc6K5
Bj/NNZrawyVrnY/kRzB30J2mzOSdBjGI9U317/gZ3QJymY0GGrQLUBXp7xYI968GnVmHJKar6Q3Z
BOh3MEhjtDGCFRLAc7o+leIizh2xYpRARpY9iU3o4CEJkTf4my+/f91MFUqpQkSSZOaXw1yU/W+c
lpGOdSZCiO2/KZGQceY0ZrEb/epSblQhxo+3hmO8t8x09RV2So1G760H7Y7+Y1M9azIYWVzOuY7T
eaaxXVeEy9gv3VDKcYD5r+JAIcoSfee8lmCYdq/2yFxVupDNBUNOCEYfx7NSHD3dUQHVieXQuBwP
PYNe0LZ/62HuyxKVbGuEbYDzC3qHYXhCNhU0CwswZPYAhGcDCvxWXgbZpO6W5mQ64Eo08x5I7zxs
LfIqt8tKFYIfkoBwBc1/OjmpgNhzZJSU+J+D+YPIMdRHAgkzXxNSRRWTXONHcH2uXF13y3wL1zAv
yPR8Tbk3DfnnVqz0OgEDTnC8BfpHKQs/Im2dfJRKcNW+Q3L64QqkpmnnXhTmaka/J2jJIE52fNp1
HIo0v3NIigO9xTTHlYihck6o7e1t4V+tvGqnXFCVqdIgi4G7l9x2GK3bw5wC2F1ZN6I2gPPapDnI
2rW2OKTXrQkKexUWkAKsqqsmF0sA131CMsKMnvWp3h2xuNgTSyGKrjWiNHeJqokPjwCjrfYOUP1x
7xeUCjmqtWivx3M63JS46FxF8AMDcwclMmRccuxlOHstuFCC7Zf+AtntuyJAf48foR1bwXy72FCE
ZQU0cml74Q/L6DLz5PwSvbu7G8uAt743B8fikZ5vmjPH3mhjnOdUNIZErZBUxiWYdlOC+TQDNt36
0UPaYTGoNAqafoi3WLOqoTGskNIydEB3kdbMWvZkBCQhYAS0awNmRshvx5enOV+mPHq8eoVBemm5
C0sqfysjac7ggj3zkB0DolGUAlMRKk0m24IuLG4JCx6J8LTtQ8HmuRwjtzrL24dWAE9OY3pHfJwB
Fh5AhfSHYIQjQyP/5U/TcsbITP9tTSICFl6uLKzUhUPZfmG8Gp0bTi1MK1QDvPjqCtnzNXGFlWpL
fqUkKfhEVUZzOHz5lI1csQtSvHMVXnnbPi7J4IQLvbm/BSlncoVvHx5BHVxKEmNHf4kgJ/+QGmyi
0oouF2Ab6o9U0rC526/ewT5Njp8GoQYA7yMXIJq0E+U5I5FXmB+fy/aSfK8/NiTSf4bkFtjP06PG
bUigQ1R0s85gFvRoXuySLL1b38O9+QqBr7FwLXWz/gdAwdyJlIh0jL+8L54aT1pwK2R9RHRv2Ot3
ji3uUm/ii4O4P7bMNec7OTMPtUJn2ZhMKzqvPn+GrFLh6SuTBbiyh/fvhY64SCiFsG51LMUXuQ/H
hbvYlPNKdkO2+TQ5wsrRLCOIVd5kDLrdL2Q7UQ4jpcP0QtH9cFOobWoCBTl6FLs0jv/hLNYJiolB
f+5yfjHWvE+N4XYka83w5wfaQf9x3xIW5X7GuR0dIQ2uWvnNivfk4bBEaQ+WNufTm087rlSS8k5y
cgm4V51eYGFLJTGb7lk2H6urg+utpwEMwBGleokVauPcZsDEb/pfp4P+iId1xPDj40+t5RJ3q+Mo
H1JpzKw6gW483ym3pCDSsdJH87iiJ7toOccjINW3HSd8O+yhQEOU6x7F8SQ+bi80weacKM3GSwNc
h0xWZYNzR39/33uzORTcyh+V42lf2pKQ5/ibfw0O74mC/e/xCFp8N/wD7HAV92kCi88iKjwGFsmf
66SaGwrCk2VLfgzobOmud0VImZQ4pHCA+at1Lfgp4KetzFaLYLKmgX/q2rRkBzNIw5/8LhjQlAoy
YnZVB6gYwuICcNDXDcJ+U/dVkUhIRFnkLKOV4QWVppjgmujvZ4IAzKxzA3ELcDZlDPeICszVpXUP
VGXiYYmzH67pwD+RlXnqzExwTAIOmNEnohQWok3XfNRsXozfbaIZr2s1RGAYiRw3oBUSou9eP1ep
FdFzVmRHKyphtleFRJA2P5J1ofwdll4522RlrpZpJ5PMyQ6SoC1w+lmlQLDdpGCeNXIewTOeBagV
O9BLKr0z1wlST4B/n6yWO5iOk9XLeyfkZwfn8L0Y+y5f72VbSgnCm/6kgdf06XlYtMI2LaxxJqvt
KaG01nQHRuSmqD9bFRAkGbmqYwNa8zXZNR2NUTVob/FkFqL49hT9eaRXvRSRgjHcpKV+px4342pe
2SoQHQHU1weaG4qiHFzM2hQEwZIEqrSawstwqP9IB9FVW1i352h79eQPHXDTHRLizMA9enoqj0pG
uP6lrcAODZzpSFiC3vEutBWTbHISjmNiwT7iTCurd3Ic9E64ytlzTpIWV0066vW0pOXwDxOESzXi
WDl6Xncdg7QlNU/hO+UUtACWeCdoO/cHHRdA0GZ9BSE7AjVQgQYAzQXNl9oKr9Yc1GX0SDOxYzTW
LuydiBvht++hzFXcQdlWi/SrZh1kvvDfcji4kKtBg8ntFGy6FbTftQbsjYzqOK8gZsOYwA6o58TN
0ttoID/7Gk94F/1EJT6hOGmU/Ny29hHV2eT/v23AXAl/trRNfTwc6EXYn9rMwiL7W6G9J/AQvs8e
FLQeTkMumpCbr3r1X4a21Iy7WVxSWmobmioxafENgFyNmzNRLHq64WedgWfz50Vpopp87P2mz+kC
+CY35X6qWas4A6DNenG6USdWi7dc914HJ90BOu2DH4bVrRj/n3M2wtvJ8kdPKnbAzvQ4dtl2Sh76
jZC0AxDRtmsNRLLGXTGNHOdyUlQ6rf5BvQzbw3NbUrPvNQntgbvZmj2L+/sxiGiUiVb6+/LyF6YG
Wgolf3H0ZZ2LsE+jVqBvSI5tk8mmC76sSRRvLXfD6gmOqohNrUAEz9Js1UGZaeJKISR6gZ2GNkA3
caN466kGx4M4ZImE/eYJTsW0Qj8MTKVcL70cmixy3shcFNgjANvPpb4cLODFG6wO7ZnEXqi2bzCk
0gUy1oWG9VWWGqel+5Le+IDva51LWbBa4GgBUw24UITPwZyqHeD4nfybArtZCBBDRDIyHudYkiXi
+1N85WugnKsWniK0YaYwFyj1YXhmAqNC0zhM1JNM8huTTglpR6zGJSTIfHoYecpCb3ZFjPQvQoxQ
ecbFTng2pyeMKJsXNCdni8lxmAlzdW04+aCYPykaLPfVj804hGbEm/gsidUKXzHLIbireJbIcD2B
5RX6de7uBg5FRPuU42qEMJMoYW4lhOe99q9JuA4GddtJJacclwwEhGIyIt6ScUpRaTQNlobAEisT
9p/BYOwIZfnc5IdV0Csnkh1RwCdeIBkTIYKjtYQDLqJU/Nr/jSdDi2sRnaHZCR9CmTnkumDX+eKw
nWl+LdZ0IufWx638AxtGIqF1g4YVdTa9uiu3ebIb99fd7U6Pfhsxi3PYhw+Wl5QIt/RrouqMtjh+
CE9hp454EvU2pmIm+N+mPWpb9YJdIZJU3wKZnbn5y18m+9KX04UaC7pgksY5UhmX2SDgL7ZX6CLk
vmaL2jfJzElTNLLpYhmVoJ4XugmkqkajmqHuHBadfbfHZSjUMTs8pK8M7y7DHSZlYLWJiCITex1o
HR3afAjxnxxjHrxCfnPLPYVsgB+CCOsLZNKHrW5leHNFALFGFCZnWVYycSmzDQY2lMKanvN6jizF
LFUlt14ucs+n4y74C4wt6RgG4yUwrLHbxFKcafRRPHC1PFFnrUDZnKzwGahufNIGtuTj1q/chmGz
+TeRgu9eRjdE8FjUAJP6pvUVCDUJoJnayq/CakFSV8miJtwsVaxoOuaCVP6HZ5zgY3Xs2oOVLYYe
61Be251PgFmrfsQwaboubKaY5oAKyAOKPW/116b1rSLzOuLkCchdnfWOe6LQTjnN3eB0gyusGrP+
rAmH15tva1y4kWywfoGtqIhvQ3YVm++WBw/s35CIsJu8utVpx8yevYypif58o24Bhmp6ySGoWpd0
odLDAZUltO971oy0FliD5hzEnOMz9wJ7e5PMxD6aknDpzQazC+hBB3IkRg16QcheJJF2vD83OVtC
zhxAI8CtXMkOpyxuuUpS/ni1dhY5QNJgaUEBvaC2FIq1fL7XBj+6nKpos4sQgWuX80YvsVZOi1D2
o5ICTIyjbBt5YTmIDISOBD9eKjqGWisTEmP1v4jM7Bk9qhdpHmT8oSuUPj5bgGgjJkOVg2hojmyM
iwSlYRHj8sAFWLJK0Jv76TgbRtNrS0o3jy/JKl1ELfwmllEPYA1oYNZeD2Cpbxm9Sl8AkzF8FfsL
NN85ix9Xlap10zqkR3crutPghMqQxmKJmnMkbm2o4njLAT9p0qCNGTcrNnBAnatXB+rCaxRXNU8C
KO5DKOQR3oz+CL/nZBRLDfS93zwc41TINBVzeRMOWXrglpb7HZ/17HaLijHMea5+TSERYzSU01qN
HYPYbj2/FnvWKOTtBiC8Fl7rWMYb1mqQ9I/Xz94lO2NdVczX8+jZB7PGknNngtF4EyVfW5TH3rVR
S/84Wq6qXGt8P/UeQqb3FPgUKKBIeh6dwb1VBCUwqkxtts8Ortc9NRSYOcBw5q43x6YQH3NrQlTu
ZvE9esGJ5U33zeycqTG1d99ZGf1xj/Qe+C5STzakaJ2QmxB4QkNDFuZamUJD+tG+MnNxUM0h8E4T
qOTBE6oHZTe4arJ7sVAEgQ4eJcdR8YpXQTBY1AxmdX9ydI0QhWCrOKrFFC/RvdYR9W+z1qZyAf+j
LU0tnuePXfgiizckoXKg+kW+C8/5P1LH1Bf/M/K4sZ/steZdaQerYCmDWjPmLLURWIU38j70R/O6
fgsUcflbMQp0wIH4C4Laku6cO57Tpzw7ra0rEZGObNsk0KXjxKe3if5IARFxdk6Pew9Diw2t9fWu
GvU7SNjYTT9EnB/Pbk45q5cJEPIBhA3ViNkBd9ezif/JASo1YWK1oG9ZdJz1o8teVCRw0E8tgCsS
m+lid1xOdIK+mt44DDHxH14ZH2i6T/uVcj6iDga7Gf952qPlkRr9zjdqa7GQBl3tN65oZq/gXU0/
y3GaA6s50iiAIWkZzlJf0AH/qEMMRfWNws7rs78uUEepp/JpWxElzKj07GaGc4bq0SBpofp4rRS/
3AFYZ8xOGyTzHhVqEe7NCFasC7/1p60YSa0PFnQOLnO1flbsbjNlMDOxRCSYJ74zafSLyiuTHgj8
Q3736jdYtHuW10KLapV5oT2ImLbvXWGhGlFpH4QwW8pYdP0HlnopI7d76jApxhGNh3K932JhW4QJ
mu6kXyQUYB3fyL08KsGPSdiV3EQWIoXPPpCozylf4L4FGuQXw5sg4/KnPjS3sWr+aQlQcdLqqeAE
LuUcLGNtrV8dzxS3nepd+VQwYVTqC64NHHO/u7rjTBihyPLZztpLOIPa6LPlIJcB7ru4cye3ZwBJ
rbTvB1ZwQNYDkkuAwPACLlYeDDzK7Wmn5IE1l/Xn668R+nAZnalfjoLTk8ehtAzqDG0PXElWwqMn
WIONzqKvctSOsYi41ZiMBMmFabolodph8KpPQZPANsp2ZbOceiXXcY5mzEozdxFmYPUT5Px6h/Fs
eDfn/SX1oi6Ha6IhhEaSAbFLQt0ZQHVmX/Nhcu7AnGoF9T/QcnvzZRTOTmpGg0ZegwLHLU5lJePL
ogxvn5EBfTgskmaEWGNtQg0/+qjx6ak5NI+GonT18X7EqMMY0XLYr3G9qsv0KC7wkK9f1lGbmdAJ
daP3NZM3+xQ/OjGI2DUm42Wt4MXw/8YJPma/eU7IsriCkgPZOdeHenqH3OMef9WYpZ+LQXGk7Z6K
AH23HgnJI7KeEU2zu9P9gs+G/pN0TfX76qCVt0DN4ONyxwqH4ukZjW+8g14v+2wcVeixK9incxtG
d7QVx7jB0VIpmyYynKEln7V6pDhvdcYQ0EiFCV77jWdpHIQVXsTLWx4gYzhfd+QevuNFCaPfkjmp
6f3Ngec5RmGwLjj3QvmD8Fy/2jjHORiYzy7Z/F/GK5Bcv2tE/k+oQHIyKsomE2adj5aLLt0Nfzuj
NGiZOLwMZWLPPbopiIbKE+6GT4L0cPgJcmi5ZK1Fgx0l7xlYRF/2xOPeysRn/SJNUc0o/hQl+Pje
d9jFdRFJ0fu1wUsjmhu40i33/VMt8hxWvt25QOLXH0aOHv4n8jWKCTGjOueha61toEfIzQeKAjWR
gT6VCLV5mxy3sndlbGixkKC3qguSwJH4fbgTASdY+oiBB2SHYlc7yWwCpiGVR4z2OJ6Y9AZY3/ty
SfS4feQWszftAg1pr5Om21Q6uAfKeQiaw5g6YCKy8hUk4ebUlJFIXrinnTPOpFizoVnSbPXGUwfv
DlnsqQB3QyPkcX+rhGNYA4Lsk6AXqYSBW3rr5kxQLl5UXCTOf9144S9lhFOg46gJ8dDabzZjFO0t
NHYPTd7SlOZsN9duxY9TwLjy4DDBnjKendEF7M8NNt+E5HlXzOZ9vzr2kx8L2uO9vogropfjYvK9
1nDXUNzEDihGqkh0+vND87I/d3k1Oz1qvpZT4Kb8rRA0CCYoBcjc0C6GYYcmOJFY4GMd+c+sHEyf
EwEf0sZPfTrs16ZVnyJ/XQHSjuR0nxPO/u6UdkjwEW1Mals29wi84lB75XM7GUwsDAjbvs3M2yaE
+ZSBSDODlHZFivo8c7sEEAX0n7+uSNAlBBculiFwQW7ThAFVSX5eX3/qvESDB3+T2ZWk1boq4g25
e+pebSFyEC2shdkDXZHtn9vtQcVTvRfIzNF02OaBhvzf2BUtLInsWE3BdIAeeQRIxe3GBEh0NMEJ
bQwzSB352NjMP1LvVV2/JClQN8CMS9XXY5POWLdm7NSyRmXE5YggqDaVZFm8FJyt0wOFN13a/xMC
JemiAR4KljZHTFQlxVxS4/KW2DNRXSwVVlqDQMiSGH8FVupl2hkIEG2o/UKqE61BYMKcpBUkZ12K
6SZTgEN3fyBnICTwnUI2Z569yxs6efzlpClBUDSbbtRfbTQhAr1yAgxxW296zWIxh5YM2lXAbYs8
KV6V+//+a5mEFWXaCCwPuGOafbFWUlxAX9oqZmu7TXQ0bjuSKbU3i11nwjE7MZsaCuZPHZbOPrGX
ShCtFqduzRuKUns2/XIMNsE64/z4fgRUgRwtGm0F6sn/UBeEn5w0H/Zcpzntbmd/UxZ28q7WA0K1
Hy+73GRt3EopUvPczdJM3XZWjtxhYifWy30vhkSl5uNLh37isjpZNDHQRJAJy3iHXKh2YQ1hL6KL
jqLRBDzP9OqzFAxbg/2WUko571Agf42SPkdWHgxLabqL46NpIQABnwEKfDKoLgO3XZNccd0Ja1bo
futv+DqIeLaw3OK7p7Oc5c7QhYtsG+Lv/aGCrNnY5vlH+MFtjBZOyubS8r/6TDns6jHYGblhzXyr
skHhnSwy9lXFR7CYs8ul6ZEE+lxq7/h8oPjxOtI9YTWpkcHEDEIcNjyn91wiIsM2B2an19PZWNqq
84Bz4vCG7yafccrfGj+lDgq2ZnXYGaC5Fyx67NTgt88c3AUKhWnGTECxPHowLVHMrbTxVDOghGRw
DiFnWKAjBjziWHtqu9OW2V0inxXoJs38CD+PNzivXb2mrz8nt5x9fy4tQP4EcQz7tXQ7HqFljMjN
acZKCAQs6rH03uULd29fBgOwkM3Kp8c+yUz2VUKxh4t3ez7497ijMeJECH6bXuBqv7iLetVOYQur
0rg8IJ/eEba2MjdAzSb3t4oV1Oh86keAUwpDgvqHd7JUIVH8ePeWmFXTKAqs20Vv+ozGlowByqtm
VN/h35anyskPXM8wElIGBGTJ/ljZdaUATFxIg5bzUnW1npfb+PgQfFOkak3DjUPQie4oXaLrvMRf
eKMPeDrmf+gVfjRogB2VNn9d/c8brX2M+hQoxcOdD0CVgop5MdKe8N+2m2S/g/CzQByQnZ10E01D
DnXOuCQGkntkmfydls8SRtFiUiY6Md8WDl0tj+lXYuGXEhESlRWpyzwDyxP12uWQR1Snl24DiZSP
zikULuNzCaZ6E1mslLEtPueYweu2OYHvf7PWVIkuKHy4mmKt07bkZoKQZ0Vm4nTqukddZ+JkDJS0
nzCsF6b7s7WAEtsyZ8Pu/4E2/HwQ3uxiBponsbNplq2vQ/Zw0Q75mPMFGOXosNHYiS27Tn17cPgF
ZW3IH0J4T1GRCY+hZ4wQWee11mxE32PM5/oVpD7aghwZce5WWLyn/TWWRu022wmIwazX1JeQrEyj
/6v4HvEYRbLPu0/xrh29WUxdqGv6gF9ojKiBOxamm7AqR6z7MzaVAd1S5IApAKKUZMZ5U1j497hU
+fR/IDI9dFB1ped3of1UpWlJIYG7id5y/4qec1a9eCxv+7v1y2ehy2Al9s2D/rvT7AUmATKocVxr
G19BOxPhANplXxWXhoHihmzWj0XCBwycCDJEDNF3QOempB9WE+WeedvmGiiqCSAbGVtcwLZJj2P2
ttiKYTK30dKqLyuChagnWiQHE9ZV5DJ6i4J9YAPYE4nbh8jGAuNzv7DcWVB4cgjoEXUnqWh+uUCV
C7P3kT7JHmJU1U4rRKfZdBaFfvcAgUDAUr+wcff5lMR6kQAuziI7g+5OAe4in7jZ3oa3Y00HbaHp
HZkLJhaZZvXcWWB7paFV7EvwFciB/Ou/cu1sxHF8FU8zB/0+o1VURfoEBWtu5DGZo6aNIO1U0du7
lg6tzIFJeYnJO2hE+kQkN9gGuqD7XIJSFejHyQjL7zM1QY9Cp34c5Gm+z2xzPslPRu+LvBltDeG7
4viXjViwJPsvHeY0XUACvRsefhj19tH/maAOiLhH2vbubadjquUP1RhLHaLV+xuccGPFbPpMy/hI
1OAGdGc0+bYxeeoPTWhlnxHoQXehHD6F/BICq7cpIpas70V7zkWtKw60HaLbLGP/GvmaDlp09bwS
drAOUtBXRqaibBm48J51tcISy55ACoiLEiDEtr48i+ad7LmMR2NbMQRbIX5fSZSLSzOcgXz8lo/2
Z1+yqh/bX7/L5BEZffhbQfUOQM3MTVE/k32N0i/1u8OitNsfeViuDzwTJlkQUNgWkaA+X+n5conH
zd7/qmyUHEGcab2bULUge7P6RfEuYydqGCSInACTMdRp8CcAn3WtMRsvjwODqsUk9o14ETaiofgr
5ZUC5prlqWiVdiQPfCC3mw+CaiaFQBmht6lPalXTzSO1v9VoghHuwR9MOM/J6ui0UTWMjYa7v+d2
MM72W6dFwlM+CKlyY7YOKWqjRd9Xora9DYW4SiHXcjQ0Rs9dsee4x7m7Kw4LWyBUGaJsvIAcSbji
UDOF871siMHpQp7Q/IMeP/hmaOx0j+LH2Rqt3HcigJfNJEgHx1CKmD+H8uvfEdI6991fVen69EIu
9Hvs11FZnIFNdMBjUNTJ8LTvNXMzuiBgcF6LbzX/6T99KeyF6HcU3J3dW02DfaPb+/1HMTFDVGJX
34VA/DoFoGoC1kH7bZnoWnwe95q3ShohtowBItDCodyF2G4UA5OdZ5PQzkOhy1baD/Q39N0CvAo6
CfoaJXEsCq/kkJyWhnq+4cajurAjazuNVTYbyYp2Zy624zMMAkY2K03Wt3mf9ILJR0Kox8ukCjn6
IVBAVjIHXLK6gCCwSfAV9rpMJk9c83tPlJgPZqb4PszJu0/hIeFg8eGsBmMr1hApzXJnEahPiAKW
OMEpvT/5W4pEEqUL8ZkIAFGf6B0HU7NmGqy7utPuwyd5Xh/cv0TxGZjq9yqGnHMiepkNBsW5xVtP
d7KV3biR5TEXIkNIbMtOE3CAP8hSnC8r0NZJfMqHIYGmmdnCIE+Rf1DvDl12iyPedKBm3AY7ba7y
QqH+OtVpSqAZyYwHFZsZomPhnbcb2yVJ//TGP9jR24Sip7tA+EQ+748tc844oKQuKpz+Wi90MF1o
7Tl46Oo+Fp+cuN1H/up/IE6XXwO6R/bmN9h4iL0EJJb6KtyUEeXx640gVsC8guE/WEEhaeKhaFpD
MdFu/qa9lc0GEDcMeBIiEUXtCfVJ++LDgsKQGipjQR6L/FMFAQAyEvnGP+e4J+1oNUzavgPTw+za
njUjSBRsnBEIzvKgx7BwnOntS+PNQdNmLetpwCuH0T9JGfpH4rMUxLmtzK4DP9NX/KauzoitYLVq
v2Orji+QuQynwBPSjd4L3DxxJBSazfvAmtAo0OLUT2Uh9dq+jDDqmMITOFOYAVjSdouOkbTRefM+
4kjyazAFYGpo96gWBfOTQ9IoYGFooNsQOBBgyLyWoeLfbPpiSojQI0R477nzXHQob/dwgQ0pPedN
mxn9IHn1vBe3U8t7/7FgMLaLzZZngHAvf8v892QD+Ir+D4WiwXYNikazVRvlfbPAOajULxKo0O1O
6nb1/TH4KwiFsUxIBNO0/kBosQ+e7+daXgDpVIGOuq212tZjxDOtwZ9rFqX5MUyR5v3KQ+v84IUq
AiMN+XtW6+jUSVxoqucpAir24ibG1SjpVB9ox4OxTkp0lHZE9r9wM4iDVJF1jO0kan7WC1TFoUIR
XTACxXRnSRlo2ltQ6xPqF2OGzsILDpnMCR62ybqj4VE2fdIR6Fi1zO+RZq+7IIvPlIGe3O/rEpZB
7F84WAjShzZE5pmsvt81x71f6vQp+YZTZm4SiEIgBv0Cl+Ys8n/fjCcPW/+HfY7OJY9sUakOaE2v
rjCTF33kOhgV2VbPs+AUvv1wKL1th957+sV380cep545bKmKiiFGC8TH7WI9WzL4PNOIu8k7UHhV
jjkaLhdne/lZRDS/resCsTznDhJ91E2vyKehPgZBW2ICaOEGd4KP1ox4oLnJz089zQlqjPdaRCEq
c7yUq3PkSdyS2fShVPffqTngbAnP5m/QI9JySoiVPH4qR7j4Q1uTCF9u6NhnUxoY5872B3P6gTzY
oQTn6uzuS/+CUbNiXQsNA588C9q9+jkNXduD50EdxIrf2Gr2zMh+wm06d3n5gAWusB/eQ1h8ILuk
T5GWvbqtcmimRk+Zzk+CuI6GWmDbpfAuo4+/HbFgJgA4z39tm60ktiH2R4ncTcbcKxTWklTmSP+4
RGigszwm6LgFRx65h6Ajx9prah/rgT6KW5HLfu0dBaJ0MM0p4LRYpMt0BOY3cmsjfcpqOu/1lUC+
mdxzk2LATN37wFwzIKPpkbGSJDA5vDkld3qDaKt5oq7DM+eaYHT2C2rwPXyszjRGV9URku8HwrUw
U2xzC31xyUeIYQLE5yY6Ckblh8IkhtpZm5eJj4Kzllok2DAxtNZeZDuf2uO+Vbt8xWLMlziw5ELM
sChDU2VpYYPxUTIEvN5xDLCJQOld9/QMDGWiEhSn2gfqGadLKAKaZjIyZkqZISJ0NzSRLn/MP9Uf
PTLp73no3Ibc5MIDq6IHdEgKq5KLsNAatBhMuKZqBdkek3L46B+rxuOKy4F+jVmQiXEkd4D3l3dN
gJIXrVFHIHur9fO8/jwmplvIjLmh/tCTSXAOD+MIhX3+r0ksIREMFzJPROghIeLJ/pGWxlgfyZaN
/6saITmarJUMlIwl9dPoTvANmBp62QYyIEIXsRvCna5afHA7EiDSKuWpMHTrIeWSVrskRRwfX9uz
kdlVeS5CIFKuWNh773b5adU/8cox8dhyxVpRufVtmRQF8J9L7TW2AECEUtRWXHbpmdFnC7MX8SFI
JJJktx2Lbn3bQwVrz3wbOu/HMx4tjE69nD7CKX4BEZiVvraE7iRgSR57FOWTjKLknpUBiDKuqk9X
b9zwiXeaId+eIWFfl9j0AeaHYgWScpl1NCRQyP3KnPuR4pMUi+Np1hoRW7s5MpIbXjqH+sMMUh+N
RF8ieeskAKDMr+8tmDW7OgaG5CVHvqbiHbyvlckBeGAw0TuA9gNMP0DTxemxhFJsHi7JKN0FWx2M
lwdu8vf1uFCHj4+K/Kirto0LV6c3Rf8Y8bmD3hA95uLUxTXty+bV/ahSWJHhgsgcNMTShCrw+uFy
kl6DHA1fIQw90RWY7uDL/+OpGlveGyFQUK2DXnFS3crdDQscPIHzTtDkrxhDOYeeQOO+Xg2VBlaG
W52j2g5rutRDl0BV1t4tBtvTYnInH2HpDpAUh1xlhLavlQkbrPhfocVN5/2R3mS0QJh95vBMzHXV
Hr4w9jkS27Xup65Mr7MZrIavpGNsdUIOlNEf2H90LcRo8cywTkuG9bsTT9jQdXzSE5Zth8FFAxxQ
B2lipjafdmlFx0XBPgTGh3PcP32TEHH63r2X6dlbJHYtbq2No9mUsmnmsIRGIAHO+zV2Viotet7O
r1trkdRfafWQqa5XYtkQHLZApMYOgV6VpJT09WCM8qAAyMS7yVaZOgo2566MwnkyOf6wGSStMKg7
gwMr2YzJdS7EalWVvxPpfblRJbwbNP9WFIaGScFS3XVei0USk5TxA47NX+MfZxjvcjtQI03NI8hc
/dzfFmKLpDBGhrfctkuQ0iJhabx3+QxmUucbQ0h2aJc5MNMiDdKDi/qiyEsHLNgehtuYaA7LLiXh
mqXySTJNrPRJnbfAur7femjCCsnbnXSfVGAXFcJjNb8nS51NOcTNFAfXI9fver1lzyVcGaAkyb1P
bardvOnOGqIOXx5LwSz/O8068ok++xjYGinP/qgFigdhDUPSiqc9MpGp9+W00B+X3hAUe6nYIM37
IFhA3X693bBT4UBusjD71qHjY/RWg3cylyKckVdv5egygDz6IyDLh1PB7jSYPE1S6Y1ghbt0ABWH
3Nl5hF0XTOJ4H8BqNMC6Z0kW2MCeetRxB1ZQT5/xQzt7VuPd1HoN1/UxkRCEBiGd/k46c/7Q1M1C
48CtdtaNgX3RgICdAIweXJhCZU2RYYXIWLWKAakVQ45uGBVXH+GzJNVfF2i/I9R7wJicnHu2xE8j
iHboWQ+PFkfiGLqzAn845oDmZWhJJL0VXF0tuIVZOKT37s+Iq3sUFtLmMFFTfbIZO+U8bdzq7vjW
OGhL9Kc1tEpCGpdxRg3gElC0xM38FOktNTVgK2aFtcESpZvN8XbLIMTqhcbmfKHSZmx26UKk49aP
vSrRjk/LAJ92fNKF+k2Cf6/qoLnbvUkHwbRVQzgTQLDU5u0UctF36dU2poiVeBQhJdHKNJI4d9Ko
HwkhukiLXlODnhKSRiA27M5AKa9f7tfuHN0y17hGShZYNB6o2s7Lu/6wTDT7FJIzxUh+A+fRJMUk
mcbQ36/gsRAW5ygntEMPmfuFUmrrOQ9QjmhcOA/pDA7unxF93FlyiQIaMybT9cCFJIU8pWPtYPa1
OyI1zUbNzJUO5y4Y+JESwqp33Z06z+c7S4tXYiv7VuSUte09MjCoIfulLJpeIaWOBux9sfSS1SU+
FyYbFeC+xkOinLygGRbA3B5TDu33POfxWShIAHPqi8V1YJvYevl67h+NLmmEYV/XFpgYMvbHi2uo
XrCYjp7LL601Izq9n6vk10RvnLHQhE9DcgRFeTWDiPinDPAg0QDRoooid5c3qW66H1zhCfe9SG0R
tJ8R4tCcuzQK+a3MPF4rgk/dbkdopk2xxaMhyMqMZd1xr0QRfFL6DfgCZU/KgDgC7B3G603Q7SVE
FnyBwhnMcvI85/F8NZgoba8SZFpktctVFz5lfkLe/tPUmif+FOKczvTySBsgfBGBeArApJ2w1rbW
72OiJyi7lwuExEVGmd/riNqLMztqrKU3sXQekZ++yk/IV5M7JtDvfTsuNHBaJRIOo7QJ2+Zu0ddz
zgVYX0EAKGpoBeT/th9SQSfINjrcFWeac32rwAhwtRy8VShfwXEIoROy0PSJfkILA6hYq9Zh7V/r
b7jGN1a6TLndUXMCkQ5cV/HtPfIo/jUAlSXmHTBI2VTjgY7YFWmHxXrYp8qA0KAsL8TktPKePYz6
567r3vrGgT37yH5rTTtLxv5ERY+KtBGCRtMRs//ciDFiL5dnQzSsJT1eW1v5J4XVyAUu/2M25aAU
JUrsC+uM54bdNmqb/Elymh018yad+NtLfe/2fc64X9Hvyx6+N9f2OXouMii4Nf6e/6sB3AwqCDxl
GAfO7o3qPgxAvwIG7zZpr7blI/GmnXGEafgHkPRFouHmbpQPPTJ5p3FF/lIY13/YTR2skRTG1ZSG
RCQAB/C/hlwEYCE2KFpu6sjdes9yjXjpbN+BJcBcJY+4SXdw4fxlZJeF/Rb33sLLsLuy7ytXFEpN
o2uRlgSfQQ0RTP8FmOGQiza/JUyVAgYs5fsN9d+uKtxp4Ct1dwJRL4/r/Jjs0kHsOh6wMwj4n3BT
1lk+paQYs/MwGhEzPzaZWUbRM5lBO8KYsrHXZ/ri2MftfbpIE3XMx1B3fnoTPyvnPlaU3dyVAnJA
nrvzRkiG/q+8OnVcmTJDnXrrt6iSlrtCyMdKWZj1i/p7a5c8IWV1qDihQw2GU6g05BTLXmOFZnuG
n+bqwMjaLNxEVByQIcosSPnVWTy5w23cSC8qc/yX3amuq5ZVJWybWIdMFNU3WBZ75PleHTFOiAVA
SYbZtBpULFP+Y8PvMhHIYx0OyU5x1Z/yo1MozaCmThU0tTJuctHCOg0e9S+3DL2U1+GUUNK+W1kp
cUMDc1NF2bTAC9gqAXWmAtHmhv2qDE+xwQIdxVF9JAL5vc9rSfFE5GPQVvW2clZrh7LR1oZhrV3G
nKNfWEDbJektgITzei5cgZ/jv9f5DM2FOnDGQ3bZzcKiqFVXYNnYaoGhvKdUZyqHTIeBsXmUqnQu
QIAuKU5jjPPUbrFgN7/Vv6a+V4EHSKtKe21Sv1KDDqlbuvoLjZnzIDALrc+QzqJ5qBDyfcXlyBNj
nwq+480yVMv/+dHeJlF/AgyQW152RnQL3kra4iZfVh+BtKtwbaeO+xttauFvp9KWKljM0HCgWqGq
gUn8pm1Cz13pqgvea9w+/ee/KyjiVQe3fOmjFs8F2jVTAPO0a1Rqfth3gB7QFYfMcnh0IkBq960O
Zux0eNeRd6irBqGm0AITdQVu9vPij8W6SSelLiO1pEz75ecYjIqVupIHGqY3dGInCTiw63p8fhuF
fKnwhDvlNxPb3PkhCoS+hD3PA6eBT6NJkzy7yOvhFKhQb23YTTJe0XWNZ4J4B2r8/nB/68tBH05f
OxUrwQv7O+Je7K3txATgGr0Gx+LUr6j6+dJRzXmoxzWYL8h5Rrxwo5NnZK/Vz3cyl8nM34GKfkaf
uVd1i/g61HYB98DEeFQOmWNtfgPyUTtNl/5c/iBD3xO/pDSbGU5nynXZnxKjzfyZizhJO4647RuJ
Lx0PUFSicWMqKM/eC0YNSatKRvrmH3vnxnKcwwV1E8QyPdhxXHFn9lZ0+2jPZKNMQTZCZDsWFAJy
U1FKKCNP0qtLNdzIsfMYjkdZwCAIOx9fPis58OPCWHGiM/gMNr77Lj5wDQCKMP2fEOIIgEWwLLLg
uoIHjhN4MqD1ch8DmwB+xA6C5359ZubAdi4ORl2GmSKSmWbBqR0g13et2X4Cac785YqZ3q9Zc5V3
CbnBAOK5ykt2MrIOwi8Tec1atIcpQQw9jldAAU5ftQZZT0GuQsEIN3tTkR2SOYis7ypdWjyZd/q5
u2XZZ+TXRqWxAIN5HimJG3alNTPgHxbCkqKaAxeQt0I8SIBs5P3ba9hT3Vh+5nDO7Snxw3oFrxdq
JNjswkPrbIiT0XEZZtHTsWfIfbsRDauv8psEPSK+vGWKmhe5z4WpBL3dzAYMXPaHrOP1601vVhz4
cEAsQvyOmKuU/FMyoQl54U/v2kKcyIBxSrWqz/JWVTJ5apHmIHmszvbiIa1Kk+na3aorHYMSnxU5
FMLQaFSDPrb/jQGquYJo1XyhcY4tV1yERyrbbpESHcbr+fd+EQiourzuls6AbEU2IEC8e+NGi1N0
P5rzJsYf/ser/He2hMDCAYPwCo8fSukYmIjh0Tb6R18Fc0zll3Rx34e9YRSlJfwPQyDgf3iLwMi7
qp/1iv8dmNgfEXH1v565jNMnQJ+aee0nkTPfGLMPKgUgDl1llq4el5E592sgLAI4WpHPhURg4+gv
R4Ji64g+TWyQApgkYjHhGar7cmM7k90RwojTlir3EdcaXYTOKVimTBHXmu6DqO0d2CMZD5SNoDwj
pbkf5cEwIPcJmbFBHgZ13YTomc1t/8Snnv+mXVvV2VLgRJkhqhivpB0pZxlM/AedW98cAS2Ztfa3
EGO3s1VGqpMlonXj4TrBYgzyKMgCG2TXt5zUcdVdktntUnA0QsM4RimKuYsiGX49/A1t96zp3mrd
buZYDObeD741aEtvfkFUdpGyVDSI+p9CHP404lEbLZuyvk9xi5ntU35P37Z4USH6WenvV+NpkJJ8
ARQbgdetVp9uUvTgIANPMnlgud0ZKpre7RFvG9ZzGwdnG97uyZmtHj7wh12XlI5PwoAnsKB+LqjE
WQTsbOFz5UrblStqZzBr7toSmErWT8pudIO1AZtB5ExtHPcqkaozCJq80ieIJast4ShJ9byLXu2K
spPA1VV8eTf6ZQGCHYQIxaNWrY0jpcMgx2dA4/prS68LMll0SRg/z8jY55oWs93pyGhhMwHcfPUs
P9W19V3Iy1IpgaXqTF+E2CTp/pSKgNt3/SwB8ySbyaLMSodKElfn7BrHseQBvDNifRrIriQqNg7c
1ewzz8LCl02LGbRsNJ5eDKFWB7/jkIiCJHO+5zy+KCldjKpvbfDn/jPsdzetVcjF/7NVqfhWB23C
pv8QrSeJZq92z/VqbcuaYZJyH4eBBm2ManCJ43Hfsve95C9RU4NlZ0Y94aw6GdxLArsfHduMbUrz
ah3HMF25o9wJJzoSMTArc+DrEnI4H+cQ7uN1gX7Cm6y0EUmZ1WIRqu52S6sveP7VdTcOGUUyn/NU
KF2INrCQJpLeBSxP/e6raxIe5RdlO0Mz8ATLruoai3630428MxqtTA0Fa7p/7CXLD7mh4gUaCl19
WRcFLjZCtV35YXRCiZYZmONllTaswAQfXNzMn49a3qZNyKcDQq9qTqzrMmwPQKI55LkWHMRoBMPb
9r8Fvn3btCBHNYj2RNNRP5ILbn6e/QsSDBOVBl0uMXXeUHFWjbEAANmgeYgF3uX871iRkBCRXGA7
lJmYaZcCtPdLj8tnvkzEYU3IwocsbqJSmv31UOAKGMZhjJUJ1fFe7c8uNmWUwfQfKoJASapujrW0
fjHsD+vKMuCjr7JBPI8rCHwaHyMq0e8h3c/18MI2dt3DArlR5P8IXnxXAICe6u837277gJ9jeS6A
0nBG1P5LPmqDG0wvPo7dN2pqKNDZXDMgoOSbOdmROu44Ja3jHyZNqgfa8eej+gc+QJKlc+dt5xCD
OYMFbqWlszkI7fFTYZwNruJDPLnvn4eMhRlWunV5NuEDdwV9PBO47k8KYDq2q/c9Tftw7cMTHBR3
TBYLcEnY41egcINOF8uBMKCQ2SKo2nsg6Prk5uJ3qV9uNFluj8rMYGPii1Fln84630xfx9sBUn0h
xyb0Z6jfST7ZjTWtk0pcU60Yxvnefa3JI6V2z8yQxOD+4PMBcaehDvX6FQhx9RDvu3EC5w1szfkQ
SVi/XaP3MNHArNner6O5aqPjtu56VVkFq9eTCHMWMApOAO3tHV84x263NbxX27keeittqp9Uxy+G
Qhfo5VTxPrsmc728WLPQR8cMDP2oE955EQOcslUHXN7Vftjzxi1Tl3/FJVc0JZ0GEADnhpYp++n1
k1MFygKQMCmDtptn4P9OpfZgVlIw4SfgsoCk4QJeB3UupNDqDb07CcOSnQryjKBtgsWim9cqw+30
nqqfE9OUW4RljRBUI00VpMJxMt2pT6SsBbmW/EF100jRl1SEJCkDiup47PeJKzNjLEwEp76jb/bd
xqAuZvyTV9sWi34CLMxfcAkqkMvM2potbL9zHf/Kzj9Wdu+/QsKa2vWFy8ta88kTFlk4XmRkLNPu
qS7L98NMHuyKh7aymOenk9pTtYFN9WsAV4+rBkQ7Fv8mDtZqN3z6cqs4nYXQn2OenRg6KxF+0zf1
L4Zsl/bQv/Xu6bXoghlAxIxaE3EtOM8Y86v61n7CsUigTbEbxRzLeaNGFtpo8gqLdwlGPXyvMuzH
ymohlndIMvVc6EKjmJ/nfl+9wv8rKBgBF5BsYr5PLDyBVJcYXaso7ILlnVYyEfscV7vYaqjPTL1y
WC2kDuKmB5OFisL8z9s+Vcpo0eXD7wzII73d+9qLX928Qw5rd+06qcRGYZ4Ir6PNIudTw0jcX0DK
2PV2mNvAnHy4ZNH36scqLJC91DAkN4ka3wUtXuXQZkEWAv2aTou3KF2DkmOaAT2WaERsINfe/x3l
XhGC/K3YwWjB6RoPHVzgmVYx04lnW3KaRvrMHPeQNj/GmoKI/C67enS6hF/Bdq+jW799GGFGTEly
a4Jx7SLWlp+01BB5vuesBUHxPFI1VWn44eaESfnv3RoNHAisESjGFP5jdhELz5PRWUMr9mmgosOx
iIqTPIc+DD+o2CXVCVeavyIf5oAHyJDTZvwkWUWf4oc7UfVra3YyG1ml+J0lLLMOXcLvTKLyakFr
5bFkAvl7t2Sx+TYO2zYdMIhrNEzfS7gcO4QYqIgnZ8uZQgDYfKhSR4lrEqDVSwKIxRJQnIiCH1u0
fdyxvVeVCXzs3hH5ZwIwY+510utP8+OrlFgB5odNdgOMmvtOl11w9dJwoYgJPzoReNzXZSautIrd
oGnm7q5hpz8QVzvdHDQOBu2NmzWE/nOBgQSiNi1a9geEDCemerxkBqKF1389t8Uidc6q3D/IKRzv
MFPmSw1AQuumrci5SkoZzmHQtHmz1bVSqlRKivZ49SizhZI2NJu9FLfQERaksrXgT/R95r/Wes2J
eDMvdwv3mJ/8FfOnM9AZCQS5UGnkWCQl2siau3X4b5m2KWXhtdPF2venJAga8qd9zuCk6AJ1uj7N
9PytKh6YPnMq8Pog2Dt0q69qwhLElrMFvpaPGwAA/VQ6tzTAwHoIMt0go5RCdVvGbB01Xor/BLTb
8vE3IIMToM7s892sr0TRkMcrZ2TS6YrMc5MRvmRd8is/1uiGurSwwB1dptOlqo7YgHwDM5vB4ORS
DICwjEoAyXc2NN05qTJvmkGTZFg7hpb6yhSPlurHAY2cbvpPhsAcybvntiru2nmZrw7Nr6zlpScn
AZ0McNMrBiMkUGYr5dgSf0Ld75cUvdX3eI2Z9OMirkaEh4b8cjMlFkpHXtq7tKTToE2qfpH2OB91
SSQmpH97vbCZ2b3Z3hrNlc/+0Qrw5FOFK6mSZC9ZoAffws4YQ9YJUE72aXVfxfzr55cF+SklKGYk
T/5y+OT1EjSHtuxi8MqNVSV++53Igu0jU81sYYUUDTpjxeExUaQbHjufePeZktyt9QJguCOW1xMB
vmWojT+i6jvgYTIm2bdbQ7RRM+8KljShQVD/KbF9YskbUZvBGSnFerHqRYKUGkZf/bLvkEFBC2Vi
cqNDxQI3rYQsaw9RRE2MtqFbWVHa0+gM0hV8TwVdCsdv5mtdtQOv+nyGeuJwx3JoJ9DN2FGR3XMF
Nuo24atu/dxrTlIOusoqyxtzndG8ZgLRk6Aak3+8kO9BJJ4KjOUIlaBOR2YgGOVoVl3VE8e8ARKQ
2E9GvbGjTiQmmmphcpflbrS5b1mXGF/XyEGgFkAXv0kWHxKwPt4anH5LvYuCVyTIcX/hUZ5UiITy
UxXEZfbjpmDtA05TifU+N17dqgOgy/zlh9n/daymCnqVGGognZi8244YdOtJqaFSq3+L3bVC5cFl
fY770ns5g5R9eSq8h6MqtDoVLErBpNkNzH+Gvajh+w4yFa7WnK0b9SzZtPLo+RRpRZSodY/15H8V
Fld9gI74yCMwoj+xZCr7JbNTacxzDjmqO91IUVd1h4Gh3RqQxfb0QcJu2cZKWU8gXpRvV/q6m5Qh
dFDmKmHF3n+V92VAm7mTohcWG9U1jh6MM2keC9xFVXZiySgbb9f3OAUGf0az36xLtlxiOm4aiqh0
Bc+/6wDTEfobTRbdeN3tKMiwfJKwomwRCEz53CNKyT4Pe2Cm6S3XaUlDAslqv8NyXhwNcokYUfyA
pM+NYCd8nsRHu5WiYlYuwyeVw8qdaioytIksyPf77EbjCoCAKO5NOd9ZQq9FQ3yHyMrRmo+YXtwK
AXdcU8ADYab96c51/SrqhHfgoM8NndBzQ1cEpXKS0ArmTgKpsdkLeouCwuntwkfqa3HBgQWczjh6
Fixfqd8RN1v3J0hAZYvVxU4q7A1o0UlNUJGlXZllLhq7hJzUFPwAh1mqVlxVhmvrrF/qRYVQeAif
rUh3avSJm+FKhVICNLbBoaLpGW7WQJ2yWrbTHKbu1Kq/tJBRHDGYWcvXRYC2CRN3e4xcqBx9fJAJ
iS3DdNUmHNhgWVIt8YhSurWO9xkrhlJyGYmsqilPy7etQPZQiT3tmuTIYPyh4suiT0i8An5RwHGj
thmWU2lS1WGYCGdmdWCHG9pMTLKkFEM7m37H2Op5EW4Fg8sevYxpgDbkJNwRAbsaPEumHRciKHoe
PeuhHivCIFEp3CQ3CxkjpMtodEr8REwQ+MzTCFdZESOY5/nAsDB8FTmrrNF2QA12ngQkoExqfIIC
dmw+V178B+l5TNi085Q/6nGoV6cGSSqWOyBPywT4G2qcf5+/pok+FaVN5KXlxYucxLpErXN9dtCQ
o3o15Ya9dvPtmDeAwwEBOkfLY2lqC3ElETPfMKwQPxviGhR9ReB/zHXKvdBLsbGTFGmQbuZmcq3d
ifVAwnJpWLfRcLqvmmeQPzCBbHN8jQ4Pkffo47GWGvp7bm3YwteCLyk0ICXi+L/D/Et111R22dIM
/8L0uxkY5jJSkdRkZADpXgHhGjhiFXFYF9GTX9yOBqtu/xKKB0HkSKaMjy21oYf53AGDSkX1icxy
S6sOHekTse/7vSLi1jLS00vnRJcnrV7S1C151rX4Gx9YCe+A6zPpNok7D6ebu48/6S+dZdOZE8iR
8dRowdzRl7ESXayBih5M4rWqdPEVKO6lEBYEJk0jCn5Aud3zseFt3ATwFGpmzK0bWIUr0Jd5wRHw
D6/mPH8CJIfl9xepb7k+gl9cjsAZd/gsc5Dr2NRUZxrBP+as4wDnt7OGxChZSrh+vbcWbY965egw
79PevNenzJKVDLfrtJdJLSy4xUXeYi67eu/6cu0G8QHbDVLJYvfA3yws0eRrVrufnPXasS4hs6Gt
sYMR1YrkmSQRROMTOPeFDA5vE/XZbPr3mxyMzocOLwcOmXZ1pREABHy3sXmkbusOsti37Hzp9y7z
5Sji/Ynw0q/GGAPuR+ghAouqMRJh0hjQy4bq6sFxXlG+nbY0IQmKsl9Fujd/tJukNFL4/Z1TnXep
md2pGSXWZCiCSnmUWsqOa4l4xY2iyhSVmBR92nTsRgApHsn+39EaTaF3ewzewIkbcsAAqWHRJKwn
/mJQ/As5SkauP0C6p7LYALbY1kRFcnRPxRjs5X0YFnqIloBFtfy66Bbwi4jILRyx3Wq/1JHJ82K3
X2Aj5UPR49x34K8QQ4K8zGPPQGgFB/IpMJtAHyulQwoJNlerI9+y3PfxCTqmsMFQjAzOn+mwlCvm
wDS3JqtezeXXNfKVuis2MbjCOWOsSgW0ao44CYYYqRhJzEsff8lGuVFc6wdy2PNyQriTRbemclRY
OdSAoJjtHeq96xfelddhjkB0ZPCq20eKZ6HeHqOkDf5ZL8ZO0bs9wGot6q5vjXLut/4jdpvmGp3J
jtU5bhp/jwILBNi8ZPR7wumSW179WF5ry/RrkOlgniMRdsRI7nxD8M4jzSViZYnMKTkaKYXlUNDt
N4L8Zrty6LNXnDBLtVjwwxSmo5g41A2Dzaswg/yb9WcxHRHNcyYy/5GfPsonY1VSKwADH1T/55lC
0f2Cr+uLEkgcyM3q62KlNzS1KIFyS12SX6BeRSe2JZfxbWbDdXFtEgBHskertIbiYDFf9KxADQka
yYyNCQtuC24FOhp3nStt5e7zFR5qQYlXXAl4KOFyMjXwN8cIKTxLowEobVv1ZnStyJ6SV2nOy8Vf
xtSllCuybbhuoA1GvYZG8JLBkzwgSIgR9bZ1RBARBVjpKnG1IbAVR8XGSOzBbYXQYUZI1tWT/9lH
CDPHs3cbtcC1e+1DVnB7SMxaMcwmiIvmPDqf2tBoHxDb0dltynuhUbFwI3VLO+54ebsrYORLbXQc
x9b83uSc0TPOjgU5KHqfKzP6tfti5PxzC3d3Wkn9neBBKYOEMIoqpXe3A7e6n2msU454d9/+ngek
Z4KwnSFsx7omGEgKYkTPl+mln6guIy7qJOWIKqEDauHw9eY0ofmqLUUtBB+wOeXk4zAwZ/Q2XEj1
4b+vgYYqcT/4LFFdBiwNNnzr63gjEq6mmW1xvrK7+VLwAEMfQpQe8h1dVuaBp5mpkPiDXwEce1lE
am5/q5BiOaO6SNYu5TTpiSeIpcXEt6ds60bTf2Ry7wIkxD7KM9cd7r6xpExAx6eKR8GuOztGnL8t
c6qHkokOCNWvZnCnj0cGlauKUQHrdmeMsc7QMcU1ejQowRpW0YakRva4fhfQC6JaeT6w+iuNZ1ji
3Ic6lAHK+ynJS2DsjWYThs9S8PCzz32FIteBSD8ze4AEeZ/WqSwluZ67Z4ie5Zuh/zcKdr3h1tiK
pBl7/b5HwBKL26HkvljxUFMt+4dcdYLPa64ppV9J3c/Gv/2msm96tj8HOHxbcNvGXvy+S58Ib70G
vdBY9vAbUrPplro1Lauhmid/RXpWAlbcWZ3zmice+wN3Q//rUuXk4PCUJ7R65FACBB/5iMBzf1N9
JWHn9uYwIAPI32a1MdVWwGlZlnpm7F0PGuBRYMorJQLyUbE2EkmpS4pSkZLLdTdrXMVn02f4YbgE
fdY50cfvXM+tx/oPV0IEN/BJYsf61CWIdQ9jPj8OEeEz1GCIiL37qqA9JdRv1BAZ30gqLuggiWm+
u/MdRL8LkZjj2BrFvCoX/vfcKAiElbLwCff8iqQT85Ro1mnOKA9Mgjrc/4bm3vDvtnLjtIxJOvPj
b6w8z3Gye8rEz7/FxM9BdhP8q7JnWINvH9Mj+8E8lqlm9LQt2YdvCz4Z+nb345x+A1AceDVPs0a9
EVdN1CnY0gh08nWvYdJ6Ku9igkZu+zE6BMlit2LUr9moUbrlSUml5tTEwt/JJ+CuoympO+Y3qu0u
BEyFp4paWw8Go3r9SWZhacebCvfM/9ZXaI+kNTYZieoBDet3b+k/CHgBrwRUSdpPqzJJt1yOSkf2
c4WVQ2vG/1iczd4J/W9V9knRDs35qCn53VHSmigRAt7+2X8JoE3uEgGFI8XiVbuJSJFWsK+SMLuh
lJm8BEP1LnidavLeG0TuPE3isw28R+S2swnPIJMTjw1XZEvj1dYP7jJiH8EpRXM6XbXbbnC9ziYM
+IVnETxFAEkWMRZOLmthxWGjD82AMBUX4/CzoNUDfbLV8OcECvFJfgAfCuspZn732Up+GSS8PJ0K
8/TQcw2OsWxLXWJTUbqgarpRf2H2gggH4tj0bmCMPGcUadk2MbzaiDQ21YgzuyyDxF/i9O2dMzRm
FlznIQE59WOJZPDdmM2sbyTrgKkdYABAYFfTszmo6XjHZzBjYgjK2clohXX56trB5SInXKE/u0T6
xtX7NuhNefynkGj2sZgi6TVYqDAAbjrQgDVdNNfFu17UFQS58VKXXgubeYWEyiToBwSh7wWZcD7Z
UK7BtVQpOhqM2ikmptSpmBf/rHW7CtYXHffqTMjjgU9a0aEVSPRkkbusaQ3eol3b5qYq9tk2y7Zv
SAtyPx2I4krX7Ag7ZfwULe7lx9Kw4GvUJcgW2R3X3sbaZ5Gt3mFglgKe19oPFxNbzdXnn8HRY6+z
Dg5NOwqVrmgHEhVMnWWaNkGqtlLUymHvklEewXqZDzMPsYQ6TMZMK6bA1OUwz3SUIfijmkmVcGE6
OzGxIKqD8k8bN4wkQKjFldiD8yGcHWOoaDioehUhqFoAAuCsCmSBCRtGXB5NNVqX2GJT47eS3AoL
XBwJ/aqsEHBz9w1zWkakXT1CaBk4iiH8DAZp2t7hWzMbV0hp5PZDbyyQ3RqOv1fwmSZ822tFkPIK
vLIeo7obYowHpld14TrvrboGlUFkGq6wPjQW+mYYJsx33NPz/VKgTCE3OKMuHMBkOrib2+IdvdQW
ue8ksxX0liKkmpD6ls/cH3anENJuw8PEVkqU3j/X1wDjJfPq/uED5PWmgSEKgcGXYLJrU5dRomq9
F6ONGWEPmJyOKb0BjfM3rhf72xHWA6C98m2kLXT09znQ24u3JAXh37heEEAn5CYYs3HlS/OkKw1g
CUxpfP1DUDXE0tJM3Ubj/ipXBpM1EFIwkE9zKSDEdn7n+q6+xyknZunBdth8v6hgsXrTf7EcNcYU
IYB8SMNajEVVMSvfQ3FAMbGEEG9AdHXyt68aYocvugRCGJ3R8nT12ebkDZzvRUg2gM9K7UwEHXB+
+A3o9NR2YmlSVe2SasBz6KUMnIRpe51hEUJcjr8pcb115ldS0imEYZXZMtxpUEJg7yhCs28Vs6VS
lw9iAAi2U/gTRwvsaCVKkuRHNbPE0anUXqDqxdO+C1++O15pvneKFrcJdoyK7MRmLn3N3PmwN7/9
S3jSl3OQq5SS3xQeKa4bsvtHVvAvHCnSh0Z7rgroUNZSGknjPY6CwsvydNvbL2ejgF0Yl6LpRw5v
QJuXh/sMgKUDvPzrM/cKJ95XIQd1lLszvZt7d0bLp6+uE/Jxs/bBDdfEfw5N2kzzySFI8i10e/34
BIM3QiOEmtGkU2oDdg3Scc5bwtXjCh/vaeVfsBIHsbcfJB+vrxng9g73967lo9NwFxNZfEOI4YOB
2dyya0MoW5RKDVCICVPdKA3e+LjI1+81ghdcOHJi4hOkMXy68qgNIF1UoTdRUsXQkzsjQ0nqCmod
M2eVOfMwgrWLB+ijwRzdshR2ycviMJmoeplvN5sCRDJhM8H+oMO6ie6B+2CqlmKF05+0EO/snWKR
IrsqV/FVL7fNE9K9epe/1m4NP7P4+hm2xLAt2FBp6bcVTnmp3vwiQQhJt4JWW/tmWOo44B5nORR8
cVstEZZTqOFxbRnhaX/h+tv8LXBDCU6R0iVZse0bBEe/X2khABi7OYCZdvmOoMt0ALALVdqaH13Y
gWY7Z7orQ6uycZkq+3JzQbQfxzxOkFqd7OqPgRAZWpWN4U9Bpf0fVeI/mCHkGc/R+PPHLLJFX2wV
/lGp/GJzrKQcWuT2dt9lXwkOkOMKEAhuKaJ02qBSvGnCpYRudpHwEwq5qfAWtrOr9CU3W8F31yab
NrVGOqni9+QEeX2FQvzXtQ6ZUMiq0kaNcpwb/e2IPVDYQVdbQ/Qbx1uekSbvL6the7mTwVABK2TN
1dMmYxaNtGsL4pWntQluRYTjLx6zp/E36Fj2F3DoUlj+kes8USvU0LcKQRFPeBZFoT4yZJP8xjbx
MEfh+bbOPjtBqlvHOU+5+GG0hxLEr5wej9xJf+dE9XbtcrN0cr2YO0tHxjscPDe481Y0m8ScpYYL
5fqPYPxeoSX/cmtr7u7dZaLLXR3ZWTYy3XO0wU5L7Bt17eISXH8pyapur4oOH2ny6pfe/FIY45ja
HNt6f2uZEgfQrxZYzhKBvOZoowi+WUndvBvFhF0NJgFsvMFbPSFJMA7+a5ucAjhB62HCXufDpsRv
XvRShjOHDcmBrAizqqDSzrQSZEgGjaBDI1h7xg/4ZT1okGbZ6I/eLbQdIPyl5QFW1+enourqouXX
HCCvIkulE0Vu9H0VI+VBAVx+EpN88hsUcirKtbGcmX9cYOU+XpfH+MSw4UlcMr/EbLwHS2q/7KoX
vwCEE/f3QYdioMsvYHfS1WzO0RW0Pwy9EH88E6B3K0M7IxKQo9vxL8m+Pv5pWcai5uq48Mr//B6U
v/EyyqatMEedd80BFD7tcxsmeNziqeEZp9YsIfW9tYYfok13ZXVUUo/NJUgh1prNcB8LQbeTmuno
UY0PAWhzVwinY1J5eDXmMwGVoc5U32mD+qyrfzJYIXQwvW/7WuYnMidc76bOqWAmlA4TR59rBWPN
dN9BpihrWzATuM2Vx/2s7gkUV/axYk6Z5FZjUF3eN/VJRDJxs8cTkhXfaXaAppucbIzufSAbZJ78
ByRuCkqdmYKKSHsOSba+EwPMbw5f1qdhFp4Ne6hpbmU7csq9A7CGZbwk+FX1TmeAt+SOMrQ95eU7
TQDJNYwBan7b44ukPdz0SqK9jvnwOeymCKYwHmlnYhzXBpTwJ9CB1ebJM1aI+r9TLllqA5VHeS3+
KSnMxNQy/Wa0QEQcnbmqblZ18NFE3Duvj8QhkKQ1JSltdSu/qF5idrw1XxcuxWBDAMcRjv3TFrOW
fCgCGG62yMYjVELxxfTig+niYMCnxI7Mw32HdDdAN6kVoxEhmARUsPmySFY7MktmYwtsDY6ob0Qp
ueGzGYqHnt0E+8dDTIIRiubks3PY59VKKYvcDAnVp8f1lFBoqfS9pbpU/7J/QQD7zsbpHAcmmI0g
ndeMtddPPBGFJmrWbmKjtC+l3L6lD94i/5nf22WiNYKgSsOUc2OVst+WY0StsUKW6mWESJ7HEEwb
UY8dWk8nVpDLYElbzrWz9nDddGZNUV3BctP1lh0ptY35dEQMtUnkCZ1k3sXrGuWYf6I9eXU/f9q2
log5h16K9B1u9Fgk5+CKfPnDeNXJbdvYQLpqExShi+tLUNfYuOitajfqEpr8Ssrkt69ROdkgNG5X
NVLzmeP+dOyyYc4HakDE+TG5wa6esoSW+opRRNiFqd/zvh2N1OFPWalaUkRu13AEIM01ewnEBOGG
JPEbbf8XlGoJiJElhH1Vzv19h48+d6KLR2f46YTZLY1Hw1zMa8G19kYqBCa9uIvX+P3PVFGCNDex
uAGubKgppl76Syx5RXfTo4mpexQ8kWJYx4BcSatvurELFOYVCnoarDk91yZi3y6+t7SQGBR/m4Pw
18IxBsABvTvMPeGdcnUUW+gixP1Ex6oHzh0HUCR61aDfSPgaPQjmLYLEoM1P5trrLSI72sPuHsWM
SBmwHQ1cJ3h3egBOfN4Vrjd6AKkEyV8Bsuga/3NmYu/n+vosi3NV9coywTuFW/XPTGZVS19k9qJV
bnIC9uK0Zw2JVOMhspalp2hizvP6MNcXFxbRQHDwboFBr36ZtdpvUinH8a6qNbKVDeENXi1G16Hj
StoevS28oaHAygX0x9Xn54cDmxzsw/E9vg0ySJVBJawmXplrU/8y/BB5bJQOsAX9MQcIKU+WURK5
NcoWuSGiDiki+L0lTwyL2MN5Zl9BqPFaymH4Ke7uRnQ2ZRkmuW9lE6gtj087OVQXng9DcJfNKtYz
GOWgv8UGxW8+iX4fyhwqIDhvfTgkQbv9sED/NlSK9KZCG69QnZBIgybZv6EKHx+NsNrNtkzZVVuF
l2tT2hbQMwdlnELmAy8PN5qu/ezBUGnULXIGR6YSJqDgAn0zC/BRT+74qRh6dp3amvBoy/2C1S8U
OGXo8TycVEDPGIwdOAPfHS+DB0bAtIQZGc3afqgLDcY8LwFBv77GBbrIXxrNKmYBOShshb9ggRa9
S/l6FXb08WDEDseB2/IAWqW4hq0TUvzTHrNVqSMN+Tb34SRfTNL5Jng5WMffD5j53dU5+IOPLytR
wqnFLqIzEtt+c1HX46d8FF5YciGF7bVzxAzd6qkpjc9Z2sXZ9bjiEFeCh47xdp1ZhQhhzPHzxaJ2
ktHUV0ddyqoIkfZzM+/rv3FpWNEBHamt8Dq9oofjjsx1ZYMCwS10iDJwX8e+F479rWQ0WdyeGluy
rC3oGcRiRYjqoOq/E0BKVSQ8vJp/xa7QUcE3HxTpq+uNf+e5kGH6G1bdfUhiFhsg9NU+lLLclY1R
Ll6+7ot3H8HPCdY/m3R84FPV90H6qdt5rflQitefDVGwAju4wo9qhPd8VYXNnUlDO/tSodgAGHja
n6lbLSEGQQJmnyUn9wYLlDSaEk1a42EsDmpE+NNeDDfd5H4hyrjvRsqMKEi11x3zLX41vMWJctDB
D04MS8ztMoNNHcXjUg5l9TyFSNmvggVt2ArTL8ab14crwIc8Xoi0t3o85nXg+9Hb29zx+1Gj+s5i
RgIcKJGM5iodwCuiIkNblC8F4clRH54NGPUmk/G7GuFqgqDgqZ+TBwi+V66xvpj4qG8FH0gaCbBy
NHvqttJtg5hilPCje8Cq6huthBhkbZQhoZzj+gOr5H+nh+ak0lUInRmbj9Fb9N1vtq2TLa83A1XY
RCxVU0Dqa3hL8SjPhyhvtpdSmddzsjlRiayY7yGZjcNuMWRb/gO2RemuEHP91mrUnJfDVpYdRhQE
XlpdM/yXQ89dPZi5Sc0p6MlkpRE2CbUDjfv0id2p8FwRX080Yvfm8msmV52F/B0Bskep9TZ26bSf
7jaMESQvtWPS5lB6F73ymwdu9qrwtoh1pkVTi5txMo/0MniNcw1U0IvsnLOgQ2dCwGcsLVYeebl9
PllGINklw/YmtJUB5WRfyhV0hGvN9yuuSNNdwxkjHyhk05LmCElcnrQUyIeQcKr3bN9wD3V6Xatr
vBdTDNaOpd+vKYR7tRas5FsPlvNx4L99oTRl8cCNRYjDSjfnApBq5CubWlWQIkxtvDfxovIENAh7
bvS9NUAC3soGb1UIMocQvZeHOon2KulVvWMR8eRek23KBAw0iE3nDiEX66tqPyhJZoFLVZb0Vk1L
wLP/Xktan3xXBIoouknsQJEhRBtpbVr2GPzT9CbfzFJ1lt3G/lwb/sBWFDHHPrdmMCAb3EDXIoiR
WiiiPexNRhtxKNvGuDaVWRRdTOKboJmkFwXs0dV+d9WoseN4in/QjHoSjPrg8gz/WYhuyRabK7Dj
orXXUDQbuvde3WhXxCHtYe2/vFkjdlNkl6esYIpPwW0P3Ox0zF+CakUnh68Jyu0Nqw062RcqxOkg
H8RGd8k05ISwcc9CrM+iJ3t6HrpIGzpH7at8JCBg1OVoEPIg0EyHEv3N5rNxYjpso8GMe2v5PnRM
NQTafmkfz+TNuvZrl/DhvxoopZMc6m9x9hEflu215fokCIHjCNXQ7wGNQmJ8OAv2CMMBrq8fxd3Q
tRXQdOJtY952Qw08u1+U4JMgFiw8cGkrtm1CFPcK7QmvtaF7VwkQzpQxnKxnMexPJR/5/TaMKEru
hAMX1t6PDYE3jNz+CKNu74xVAyv4HwkpNDcA37EgJNhMm0bSW+ZqwbE5lU/sKLvSmZANybJs5jIQ
hBoln96ow/9emBbb9gNH30ebrqFhTxxxjt1OIYObJU137YvmkPT621Z6DNosaumaEatWvDR0K/+F
Yx7QBcRvcTT2sclcvB1l0vF9d0gZlta4y6x3vmugqNXLez6LvqzkDZ0OiKjvs4taT/grPmjFbb1n
jabDpvqWTNkmfWa8C91HLOBd0vvk5JDPfh/8WRVtBVjx02VvsCQjc8aMUO1T2CkicpRra2Ve6Dou
CUwzVhXBhkFJGVHH9892ZCbtX+GhLc4DUlM0NsO0/IF0OuQHqC+AWpaHwCDkO3U3rgjOwGUNQoba
jMZm3/W3IPGeK1SayfV6qRgN4Q/o/qFj+sJhmidJXBZZAGyeBTpE7D2Bnfireur9IZlKNluTP0Lk
p2iXbitPdr4zooJw3Xl76hmttvVePC1uN4UvI9QYorqkPXptCPUzPAJGpVP/BeBCQ9mv2W6EWVaT
Yi064uWznK9b2fLtb2u+qcjPsaFvlzKFwE7tCL1T0Vvn/KCzhTePoqqWOw/P4mbdRVwKezYOhTr9
SrdMVytX50aP13jJJc+HVhXoytAPBX3hyvqbBRbwkFmujJtD8wdhRLf5mOivOMcVXoonzdyMk3RM
4ZBEstN9w9YcWkbkHTmwk83+7CumpZp3sv1GAO0K1n3JhO7YxoDvQiAvs+rSVhG8R+KJWyk+6eoL
sNaIfNOpUxn+Ga/KBrKD7klvHaavm1UTWvSFCgoTF5mLpaVsSzaCXTXH0VT/WLcr9QRZmTZJtekm
c7Agzmpcgh16Nk5II0pTUDbpeLLy1IB4r7ZIyBh82Tu3t8WEcSIvkuHyFA/KtiObDBSWg8APygmd
YaZFp64r4zGnzpIJas1RXz5ujgvrEjTNVcbmYWBcsoKkznwPpSW3/eDZjP2WOf0/wJYd3uSzkiXs
TaWINl/XzwSSaQUYbfea7d7enBS8n5nyHjEIvSaJv9iFlJ3luTx0AXm4Ej8qCzzEf64p/91+ndqB
84PCpu0xG4R9jJ+WAsswdyrK2lVpjSmko+8fvEsG9AAjLwPhT8avgKUb8QKSR4F9VnjBrOI4C01I
6jvCmXgScB9+LxJSD7k7qcEjTIWCK1PeYvEqKY75uAD15EUZcj+XL6/YrPddKrDJO5wDxU13U9//
EHBQyhV8SG/Ye73oEz87LEm63Mca5sJdi+x4MS9a4aol2dcf2Jw5mDR0ZKHJk49SZGCL42Grn0z3
OozYvc5LO+fhVYbi2TYb0qPXuwKnIDJsUKpnRWL0Ta1WeyTWcjs1RJmTO7l5JujiV3kav6VaDQ0E
PxoAfDUxcKZqWnTABa7cq+L1G1wYp0G3Fdqdh3z2aKno4zFW3S3iJmSO+yIIHbewmmvfkw/P2Wd8
d6c32/DPluqJXPQ1aWF5EpV0nPKo5bgl0WZ14hMyUbOsPgl1e2e65/QQsEZ2sWhaBVMdowo6kX+c
zfNlQzbR36NvsjB2Def59ucT8se261Om8NHZPEykdooyxzL7HUN4uXalo7CLPLQDOTK/CWLEsdDo
CMxWd92ln8MCVFWpMBzjOpPt144blGhc8a20Ot+NIX1qbWTu+bWpjnxnS1VAutkZod9M7aG8sA58
jT650XXX/k4dMjI93bWKpTYMZ4lmNiWTHLTLv0jEXFpBM2sOWmgpav5x4mIi2DpJ1PTukvV05lE2
O/Sg/0TfqfKTp+fkOrZjMcUHgcqSYXq6PRbPDlMFc5j3TopEQ2biWMDOP6N+yfC0cmnUxcXdPxQS
gE7aJYX5uF0Ou9CaIUQBZA7atif0Poa7P7ub5Msm9Xm7VHum4oDHPAuFvO3pVKrEGXDG2Geu84Hb
Z6A2HCKKpONPUyqQFKBKINajm742I4uEP5iZ4Om7rwdVMiOkJk9qa40plRywCQqf8t/QZ/yosI1G
kmUnI/wezbxC5DlXtQbuy0ZaPrB323rhgLOUB4Ahke6KltmsvF6AauOkDGuD7Jydw00YLWVR64pR
1MTvC5Qw2UfIgbkG/olAG6LRMWoTmPOsOzeUQkNvqjKeB/ldDoD9pHwpvljRfz2Lfxm8UiOPwTR6
1UIlitLkLcqd/InUwDgr4RtAwj8wbgNYfnj6z7AHkwqOKVKIFnJyzmE4yu6vVyAOXmGw3Y8ebZH4
KHNbO2BO87iYb5C53MkKBIhfvO8F46VhjCfkJ4MmPFBlw7gzb40AzjrmR1JzioDqs++XzFRrpxqS
sG7AVFLfkNRO2Ayo0KzvvXcjvwx/ZmlOp/Ou/R9pTU9hZISBljhlvpm4nHQcF4Grba1R9Uq4UQBo
z7bD1cammrOA4ubEQ6viQfZBfoQtetZLLkE4DI2QFN00y4taSigQykpUe680qlQARHM095VVs+9J
/qYHw4MffbHiq5pMn/XTOQpFUF/6dZLpXB3PYvV5tr89axFLUjnihQhgmoULtUazMpTI6pNsDZyi
nvaYjzQCgv3kbkXDiGAZdbr1tMiQQJVb8wKSDhm+uHnDWVCB34THHvham1UoAVMsg4rxSYyfLYql
ypuLX+XxLqLIqT2cscIdiRHoIYsjG4xdP2j0yMevGp0/ub0cubS7GON3Jp/Z2pXH6AyhUJguepwg
f7Rfv8mLBiJjC4VF5rRcT+BpnHi0cCqV8jJoAA5wP55tvUqM8KlotzuVkhDzP3KgZDlWM2L6relu
Vp7ko30IAo4f4lhx5sZTn7f+8R1LheotTnGiY8RnwxY3C92EpyDdeC4sW13jp9h+M91l6XtyEcBw
Tggx58+dAqqUEeK76Biw1uCC9Vb0nWqrfhLiFLez8JrYJE25QmqLuU9TQhdCLPXMv37w0CloUn62
jttU3XzMWDh8LV/TrjS6it+TVDT4NUPjvkIXeKNPLTtyLaHwIvN1U5g1jw5HDzvPuFqMe2ZbQGHp
rwQBlYeVsn9YOmhsm/ZUnBi1cSF6AJtOPZcigl6f/Qwn1cfMAOX0MAx39TorsdckYO44f0WWst14
g+ambiQ/jy9jhdjwPaFMWT1J6nAaeaJitONwSsixqEq2lDYp6iwZb8KaTBNJ/JfAsX30JRKiqZw+
FUMqEPICfBI8Op01jVhfP9m6reNeXybW3gH6aI72K0D2szUgLGhBRTyaSYRqzPTSOXThh1vTd4iB
hHqQbNL38VX4NS3N7XKvqTK1pU8/mjdrwFjifhK3o7O3/kRNroS4QXhXos5ZP2DXQMoB054uwLHY
ucuPy+vwdE28fmdgszmkJEFgV2LU6C+qxm5lVzQNLewukXuSqfpjQ1tgZvT9SroPT2hmKg2rVjRb
P3kLDLhekH8e8F0RGshSWN8asfU+CiwxifHOXuDQhfHCs537yDDtum0TtRz9qJVe2t9Irhw/11mI
6+j1Lw0HG9hTrF5SWR6q2he3osicUW8KY8rMTetWx/LRXq5ArO4AademNY4Rn4mDJImA8oNXk35L
jnW9tNq9WQKSqhd/FvrtrDidgpCA1LhIRDlhDjSMw8ukAkDYHWZYoJYYXeYOFiFy0F/4jLB3MWgz
B3vL7/gnSxJQUNYKLxaX3YewkGMfLUY/N9ALyLPWGm0zBOD5oMrwrcg81mdH5USfPAfOavQnq478
zLf++6G7/tKFBNnn3sG8IS1bKfJ1M3kf8SfTCP66cIbeqG6t5tyVQBkO1IT7xKg2Es9KxTiPj+Fp
ga2g0JXtxkqDACWsBmJFCvCIIsGZz3T3vinSRVAiGaSxd0VypNmolL9SRQZKywja1P84lYj5Yg8s
2YCYMOGD1Yrvf8Or9EKgcLQLCDlOVQM0ggHGIvglF3lQ3AjfJTW+pYgcbm2t9B4aySmhsx6Lb8lx
mOIbG96lxFOnVkOd3VnW8ElCo56FrFpNh1ToLA4wCTjPecZGQLfaAu4Isw1twYkdO4zS9/ruiQ0L
zcw7JqIG3XL/EPWDvJwyYR9DYKCe2JnK1AgFjssM1qLFQUPX05M2uCNqbJfxbhuUyDoCEatlOI3C
nd2DwzqMvczghUDDfLSJ43BFLWqqTfCWbBXBYyUC/yI7JteIu6E5b+g2UgLSZhfJgRRB2ug5cT22
Do1p/gnnob2y2pxaUpXEycjhtBpSVJP4KIHHB7tCTBaJtd8GuiRmT07LT2G8UVCPA1lQ9WQ57RIO
SDY6+PTxSIuquZ/U4d/dSPP7Cs8yHfizehmdcdJ8y4qoX4lBAaCL34jOBKKXb0E+TFfCtZ6nw9H/
kztIXFJiQBpxsRYGAlmOIcWbIYQ540hYsl2AikAYDK5CNYD1nM++ZuUAlzZpBjEgKtN2Cralj2ry
rtwtX+BI9jnG/7XGLfKLqAZ/s/D4RdsEwF3xXu/8qGWml2J2jZYHbjCpivqh3ocyTVzxgB8tSyrl
NjgGDDJU/oi+183NWiuqetQ8qGwPcbuhgdZ7sq0JN+oAe9MjFhYZ8msNTl9JA1vFmxKdF7oRINqE
S4Xgr0KzlSmGdQl6HsPfhpFPV4M9Oa1TNVSqsrB2y2vZfkUfIYObBVrv67woyvymkIIO7iJl4JGH
NqNj/YSPFbfoZpSpmcUer0K8dYZ7q+Jg/xtKJYzQq1FVlJrKtYwYy7eXRZ7ABgZ4ZS6YDz32gUpR
h4CC66tv63MYdrKPlHiUnrHujovVK0LxKViPqYirrCIDGwLrVDQGrnFdFVV8sjMGd0sLWkmf6GYG
DZwE0BkpOMeBJbtGmhBnO/vZ02QJC/3aipyRlqFSr856f9c+I2ZniqspGqpv6ZKM6vcfOLeOeowg
kLps4MWCEa4mOPBoqKLWncxm93GVqOXe0Y8x9wEh4YsPVgad34pkcIw/5W8vP36NrmcccBd5AXZ7
YwV/UCVZeJnM/gNmCtuGCM2JuwGmDOGCSWYevkoY4u4MJRtv/9IVqvP9EnJLQ+xai8tGhrpZbaoA
3TbcJ/K4KXh+QMarbvHdL4jpNSmT5DwgFmuGL+Qq9lGHZSh4k6Mkev9AsFRB4jQEH37fNr+Hamj0
rS/cCXNvxzmE0Q0VEYdpfjv9083sssHNPWZS7l1rB6E0F0/EkDMUG7QAhm9ar8BV/YK9Jfu79t0g
BsNMYdkYZLKeUyUqfOzUKa9nY5JEkDlsesK/qwDWzbjp0eaLiSZ6MT2EvM63MMKZx8IlhsLMkzSI
4Ar2E0aiv/C+3zIUB8LLmqDrM6ISh5vfE97DLc0uh0SPExyVy8Pt7IjwNgLY2PkjQSPJ7nbyT8Fl
KTE1uO39NY5XdK7RPpG2k+zSmYu54rnu2K1W0l7lrIDKPkmz1UrNbQq9cLJ0CqD4zDW/4JYa1F8/
B9bCzNk7iAsF8axQ3b8PvVp1pcaj0tS0w7jDnHd5T0hU3ssljexiadzTiTvcr2DgQLqqP/WJzZ0J
qy0GJvB2x2CDHOICHasVOIF78YCs0gsNpjwErDb3uO7ntwsN5XlFRHpzrTytBv17uCBc8bzXQyer
fnj50SRflQwVuoiXDUrzsJVD2aloSxRWg2rU5XMLZBS94I7acNAhiEtxMtp2HDeAEEmSyjROZW4A
x048fbcMd3WQedHhbNXr3iZMLmoz5JpOFXmSmeb2rzLLsNNjKWoOkv72AMZeHVivLnj76srqLtlT
BF0ZnLMcPSvU9fg08zRn8BPy/BbxtIlM/adqJq0XzwXJmoJQqjjs1dqZJipTw6mXkqrbQHMByS57
+hOafu0UZO4c/jNVTPbnOe1wQ1z8a4kato9T0K2VeSkl6CsGmulAArZTNo5gZUT+sLVpYqU6Q0DZ
igwa7Oe64P1mgjXCnAsP5gOxCaXSS4pIJQ+fFk02e9xNZKwoGSoWGHwkFz+RSmL7l16yMYCM/sNY
gqg6/gELwigKwsryjp3IdZUa1+xdT/Sm5jsoR56RAdJsXq10Wjh3dWN+UPeR3wwqtYe+2IMZqKxt
pAIsituvBNkn7fbjBdwuF8vBpGCQFBof9Trqnjm/riN95W4v6hv2KVt38PUkSxZZyMvLdDIatxAg
OXH3ze5cxmqZRob0uoXH5WY+luLYgP5Of4w1/mkiGhZi0sLprpmS2cdbHeDQZ49fcWvoMphhQjdb
BcmMQBYEQcgzevJgLtS0JbMNTphHbQHQVEVRa0cBYRJPqcTLogR3TxFGmBtyHcry+w/8x4aPmGOu
LzAeEXD1rkppo0VEi63tgKUzX24ctyH1mwr3w7zd2vwUFCjzF+9KdNDj3bZsn//LZDK+Hi+E/X2i
x2HzumyhwdXu7eL5tjZLC3p4QXglMOaWeA2/o6+PacvvxvIHtgHHsqCBNlYKDwAL4WjTJ4eK6ktM
FSNzqsYCsvqZ99YjWhGwAewI2jpo6ngq9OovSoeoUU4bkqzz1peI0uQMFpLok2tuhrIO4epYBgd8
+v80xesn0+xD5GxDUMyDOpxkIglCa4uAkUjSNJN5CUpe7mmIHFc9SDSlcoA2elPlaCAVUsH9GExi
MJ10Y+hoV+Ijcs1wFWiLCimnzgIgFmWqYG2ypy98ozxL/GRiyrKXYl97datcIdcZzOlj32tnvdzG
48w1dKUmOMoPsBLN/OEyDYVMp+SLCcg8Zg1cg1AbMM9eR0Eno8tiR/aGt3Z7xPPWCcvka8s+76mG
/njgPIJ29LdHL6JFps/my04x5ZDaksYW9PjRu6ixpV6W4OyBwAzCXIQTajLphaQaXmnf95DhyUj1
19/fNPNzrOS6xwkr2lmByHNM2WVbBdIOphuU0P630ZP1KUjJD0kTr8zcALXcxlCVN5WGyNiuKFSj
7A0XBOi8CrTn0064DpZF2Bk9HI1SjWTK12EZmAFfwM91yPIMhCPidW0E7M27EsY/m8D5fJMOzXwJ
vtmntsg+ZNPiD4caHESvK9l93QSCWKW9829zwWbs8eBpWwwPcUe5eMmjKom4fSQ5e93SOzuErcwL
oBOuzTayuRFoOyal9X5caxkwkRxqjc3cg4vNqiKnGDkWFgo2pKTjYwO9Eec/1RYiG9TU+8UHhVqs
hmMGjnZMbYuWJs6FbAOczR52ZmIiLLuV8BBZ31WagehtgdX1RMB737rbGej+u1mkynE7boJ9Yk7a
yAE6etrZS1cDWmP0Y1YS5TQJtNWQGF2GlrPEi8+CPOwxh3xkvW6K7GMpVZ26bpiChJPXfW7E2V5V
0soei70nbXsibtVYnYg2Yx/zImyaZWLnFNQLRAEJBwgnf3qUsPTdHOrCeCDXFucGu8ixl6Xteoq+
F4jJa6Wu6IpFyUsT+Zdi0QC8v/BimW0RFg2/Gkjs23pqJeW4Y8NRlO3lQdnAkPPN5eyZHUAuC72J
ZtGI/8ha2SFagEVddVzJTvLhBV0IbJIRhqJTH7G8s4iw71W+DFGBH3oyEjeHCR1oh/9obYmn+KNC
gcWC3jZNM+I+7JyFqSIy77LghhUrmZgBmjSogdZOLIUCYI/mvRRdr8d5b6pv9CAubiq5wfeLzyM9
ZByeI4V8gziiKG1DDeysxZ/gH6ZiSgNbj/MT6kpQoDUaUmgM50tLkgI8eRrCkquRE+DEx9A2qjhE
lq87Wyj/XhZrN5LV91UgH5Mkp06/X8zkbnt8ZfXEZDlHJLWjx93WS9IkI8GFhCbCziiMtSpUQMgo
u8G+eNMPI9HSir66ZOflGsRGycE8ueUafnAQdx2cUbgI+T3fEDfJXZm8Vnv+2TLHbTKG7Qr0792Q
oonl3aPQRPvoE9mWBdimuP9Mi3lM98gqdzFapjwboTrUl9JfLB9N91qhDHElgw7fOZmFljXaaHkN
1KkHIFXcjIcVhtegXLduvR8Vy3zE734/EFf6SuT8qa6V20z/EHYBW+htXPtZwZsNWZaUoA8/S3gR
mRdWbLLzVAxHyLyw43eROol3IG5L0m3L/t/MQuvrv24KRZ3+caip4FFWvoypwZ4gH4+DnU+dh7Mn
8a4kAYfqfoh8qLZuBRwP5wE5RcQenSJCcVDK//MdRSIYo7Q+oQvJTiIffxJXQ46GwGHqjlNkmK4w
xCafPXzouCErvdXrg7g3baCYmpKVdHXPq10FRUXlV2pIPhC7UMnurMIKblRukAvafGUyPQSAZQ+s
7EdqCS4GwzMUsdNIqWdh0fGCAFhw+m40CJvzjvgOR/41IKqV5Z/GbTniDv6yJze1oXmrjvxLW7Yz
t16fkAwATbC/uvLUXifqG2nOhficNIoWOSnRZ7xtj8JpfEqHktOIuA5sW2fj/l2RHVZ8tpyWz9xd
mYznOz93+/lJEEQhwCx0CXzeGEtBOfysdh47pjYQCRTTAaK+rAYiMDpveHzZ05OhLIAADX+dlBMb
TAXVH1+pv9WBUHCtazhfQu+EB98zOB5w5532a2yGeoWNwFutrymJzOGlnJqSpsjAh8d17slpCt7v
K0pbcqgB2ls2jDwXwY29WhU4+DpdjlQ0+NcMItqZXCmA4loCgtcrL8i/XW/W5UhZia+wcW1WMOWa
dkCSN7a0ZtsGaWzZveK5l+kodtPM1K8XHD8LqMqdXf0p6psSgPvlyMm0IfKFNiaHA/XTFOXaW3kz
wCPcaaX8Z8fiC7bQAHRs9ra5guFrcO9KADFW1ExdkJirDoYi4x0NQb8hkwGpxzCBqA642kYLU9fH
zZsPSKdcWTRxKxSXNfhqU2ZfK7X9fV4M/SC8lz7R4FJmHEQ1biInLIlwoCR6elj9favgpwTBSzmH
kyN5IvRiH4f4G5REFC7WnyfoYC+/Yj0xwM+13dWK4gFDmhATcUAVPgZKVwJW50agmw+ksJJUwZat
6zJQWX7QZrMwoQzNSd3e/tZw+XAF8PzmG4jec/SjXkZLAnXXFfsDa0XdapA8VVkPkZI7Dm033fbt
21LJSSECxES3sS02QUHRuCH08ocRjwX2I4wrBu8ROPpy/Hj7WvXk/ibCkf2suWsrQZtUreU1tNXO
s2GIQDwBgzMxuDX0ExhOHjCnlcKlGihUbADe5PSQc3nnPuQeMbt3ZF4agWFxj1OtlQoghFoa0K00
XkYEaIcvJUyYJKEgSyEwZ1g+d6s3SjMlgrAqwxQdkJmfB/Xjmz1WD6vFQMKlEh+NESqn5kwt3CgV
E1VBnRRBz6WCk+cnfUBwsxFHjDOA9qeLxFkVHnZPPFKo8Vxn3QH/XdnzaJ0W+73vWsIenqzBC7EN
avCuYT/FwQl/KsaYaQKCOB6yBV0DOWFiv2nAhjnpgttlAt94ELftw3YDSPo3qa5eX5pbsh06xMH+
bfK5zcVrYm7OaJs/OA3HzXKP4hdxCV4ZTvKzfHGRN8IojDINfs6MwRmfoAy33ikjpPTjTra2Cr3T
vUpLLfr1T9umSyVrvwnYfnmQCHUe6pWo1xs4SpwUTwlEeiMep37dSUeyXKRK7NBY8KzMpaitMum9
/bUPhdkoQFyj0iB6F4DibUlI5mFdH9OFt7qSUxo/XBCL376UceeFszOuZqxQmKpubDD61C6JWq0z
aigQ5txaxl0SMWOqJ1OGh9Z+/nPGvDhhkP3jKMhahuMhHdw9WDu23COzoniCWywRIu5HPVDum7h+
atkhCRRt9GHl7ujIZ6MepSwtyMlFd7wc76J0e2EgtlyIgIyS6nzHJ2upcB+PZK3K25DYmafoeJ/i
I8dPp7UrXqSSFJ/IrT6cuhaLGjhfzhTepEhjhXOj++FbpDSFUAuasjIWytfKFCW9cOq5eiq4A9ln
JXOXAKK9AwXR4Wrh8lsmqMQj1th/mwBINDwfGvvJxmakxbPlBFlf4J/A4bC40itcMVDxiU9ihh5i
e63GJX5oaVEvjvJIoZd3Xc55dePWlU3SdssNWHx8CE971nB3mAwYpbm9d8v2DjpMykPdstkw49eE
+eZbUpCsH7NA+KEtmea/PPyvFoTaTH4u2ek9gEqjcDjr1AzNKwckr93MVCSSxXy1HjB5tmp9rZiw
/SDpibk6Li+F3d3/LvOLV+5SwrbfKicRc+VHCwEPI+P+ZJJhfHkgdZY6gpM1PU4or9zbRfNQ+FuC
ox5RVxmJd/z69XER68Ht5wc0Fv9hlMJuXdOIuYnwr4ke9r/NgiMzb+rBJWhE5TVnBYrSVuLwOYtM
+wtUuYn4ZmjNVpjPJrcxm8++5ZKMp6m3cjelluTI5ojuyO5C4zBQxkskzLYGXoCYKYYknBm0Kea8
pQdbTfLHnqZ4NNhL6YlQ+1WkGtyQt7LxG5nf3FxKraJqzHpINBoy97tUa274y8dYbb7BsrcJRt7D
l7OCTk+iJZ2axnEzmrC/trvmAxYmek8iWdPh9JeWPL/KOcGE4EBY5oZcHeY1fRstGpkVGSukJhon
+Zb1/etiUlV1eGSsKoKToJNXStg83Fx+dxXIVVcWfSikDthX5AGNwox1bzOfn9cb0suX+FhxA241
rDG1KGGkfcMwTZUMuxRlRwyN5NbN+djT/cRPk3DTk61jGYufkAgP3EeaLqr8+Y8wvKve3HxHRqwE
ORsGg1me/CNLIDnXjbqZLFFKgU8Vl8ktqsQppc7ovXBGHrnmQOQT19BEfLNXJskgfhyoM+xUVdF/
8D31JcZWZLqQtC7+1g+ZjVjck8qD4kqNLhy8XA+wtW2uV6dvCgociCK6kiQW3Jm1BJ5j0qBNiiEx
An09xHQiHJm+CD8lvEzrUx4tzdd/qb4+XtmmBZ1PKXfTpK/07+k2/Aekx4sE6B7DqnGwL1Hxx6zg
JlyJ0/SxHryR2vpDkNAh3xACJIX1cFpLgoMLRcnnGCa6rbzcpDd9ISxL4gT987BUJBWivq2cfzGL
QCX6a+46wwjTmk+it2/j+j3uwphFpnIeXxfXYXR4MpGgvDqhR27bdDDzitcAAaYotyX6MfEpvDW7
nETIlzBjb7DOMncIJb5vJlMsrbh9I5Q81oKRJsuvzFCaOYWPdjEx58CWLrjcljySsZCP7YKSiVvm
wLg/kTUMRX5kg3xTOvrmRm6GLA7SawiyRiHw82hD3F8VMWHxiFLAhNIBHGFUSTYO2+qqRHwvxLDp
MBphx/E+b8bbr1++uUJ0EEoCSJwCpWU5ZQ3vFv1nXtZvEqMXkvGx8FTNFglSoJTRE5Q+YR02haZq
E8CCMpxr7Ik52UeO2i9eCT8funbFOg+fY97cQ1Ty1Ev9h0hBAmjh+v4V5N/SvpBIDAdylsBxt7ZC
A6cCRJ/dgFF77sd4kAiyL0GS8dTZ/Nxh41YCSHaOkfHFHow3ffb3t20k1K/3ljKpEh14mJj3/I3K
6c1z1fQ2JuBOzNY+OJh4QgWjHB/MS6mh6XTXYV00WPNV4s+5vpBu8qH8q7UN6y/lyNQ9H/6nQ483
QJ07j+3MiPkGLpRv2eunPmMxgFLzCNawRo3OCOnzPO8IgpbwKXYuXZUcmhty4pGqXJ+QPRKlpTRa
aVGVNMrUaqXCyW37LhpD3hqsTQOrdKC0/395uGAIci2h2ktmTjJJKbnei89YYzK2lKWv99vvExd1
l2xRl5iytCZfUuLFhW1NHNfmt19pRLlbQSUb5aGHot3uP2QHW47wAZWwQNpl1ESVS6hXn1xtvi0T
iGRuDIUkWmEqdWbcnWhPc+fXTSoj2APUi2vvHPOCHUmSQ23DRwifOMF/kfxRT78jYYdINi07CRFH
ygNSx+VgodqDl8JHB/Wc2GFNRo+PKz5Ss78/6zhvobJmsHsh0B41ZGrDogqWsGSbST2VyDoNMWwm
DofwsTNXyTEDcUhX2g/3ZQhpC3ySTNswg6vXiCqjifBgyONP/KG2FFIDKLjiL/iMpDNRXm/jGjpy
W41hVXsSIJ7xUzqdfBhhyTDb+GMF4VaZaWUqVdIPKdloufnkSHc4NoigoL+HdoIFlf/P4YuVx5hM
88tItuTBLlgxMgE95H+Q5DZhSo24f0jo9eak2RGdnzDbmDmSeTCHJUaMEcp2HJ+0v54kc/P6irii
Aell56uIn+mROaqi8ttd9tp4UR9KBbhQG+mpHl7gMFAoPd/r8opgZM9PmQWwQxq4lNvrt7O/6nOC
AvgAZRIoIMmWXlRGwJkVvi0osmmLmYrHdIuric6yjccIyR9OFXTMM461/e/sBXxqgrea5nfNKuZO
u11+HyVfypkvd//99TMT5GIJEEz8cQR1mhNokjPAll/YgCt9YhsZ1k04qrAe+08Dv/FosUWh6FBc
6aFWZ6IRNa5V9Tt+K/ASaa2soSZhqJdjt6O9ZBPXx2otZMGRdM9/cUv+4vJDZhH8jBB5/lIp1AQ3
d0Uon4EQw+7fspxQpxSdcNH6kvDHHrmmUqzBmrafyPkbe5LPm6TsL+64z/coPKnVn3/YFLZTM1OY
h834mrhkVPzDZ+UQJgFXcEZzXZXHXFD7d2teebyjlU9Ba8NMgQRO23js/+frQ0PN6VI+90WpfEJA
O6OtWsONY2g2zOT00OjZRzIb8p/U17YpiRtr5ZrEHLD7mnp61JQVwkpLoYU+VitBw7zoJABBJj0F
m30SE4GXGEJFrInkQXXTnp1m+31yD5I/NHRbmeBpXY7AqDhziNyVcWAYUjvpOiZ4xgGlAUSTEhOl
xo2yDV9RhaiOxW5X9cZsiZuDqF9WOR4FGPTaqsXPh3OtN4WObUqvwoOJaQ5/dQxHpFYybpKTtCQC
7ZQ5EG/CIV6nxQxlfg+fNlge7fIwZM66icGGD+aucPkDPfLsM2mXl6KcRaM7nE+9TAFESyEguJtR
40vbgaDHqDScCBimpe2GuRTcp720KAkBGJSiLhGwhckVIqAu+0sg7WamFdyhnWvZMjJjIOcvSUoO
h23dn9C69+Yb9TtldlAjqQ9eXuqNLEspoyaYdVww14vJ/1HKBPVu5+Za1IRWcNaRknnZbQ8INn+Y
cj7LOLuoBxwEohi87KkB+gD4v+2i6ThHA9CfM+Yj7iZxEMZtjc6cVzVhNHsaLhdFa1Ih0FiRuIAY
MhfQCc3BwjKIx8BKn/w7JjvFQDAmoh2fhI8L96hSF/k+fqgjjWuVaoLbdt/Ot008VSRQJD9Trdcq
zalE37upo3JOgqJEOWpF3+AYw2Y7vM0IiEnMX8oDth17OMQ8nWWxH7AuKkhVzV8SbWGfMYIbcwF0
gtBIyFTBuCnVZ183UMuOaa/+EoH4wWB79ulraBOVOBRM1kk+Ck9oZ1W9DmTXuk8C9+oOSoFqDZ4F
m7ZAjpP9HRuypSs255Y8LyLGMOCCoPC8WBVPzAKssdxI4bW7T7yvwiTtNwQ+m3vb7mrCsGQ9b/BH
tkPZmuKsL+JX0kUYa67/igtkyLfIsamnPu6lIyb4/kiApZJXPzB8xTFBs+FOTp+MDvnkw9LAGRZ7
+9F51ThLR9fCxdAx8HwDpNd9Ut5iJVuN1seqH+R6LUuTKsoDAbPDTLhhDE+kc/zmEPLdtvjc/r6/
Lm+rS8nNrQdFJeweL7SpaEwXXs2HXxQFyNrfE0w87sjnZiMPi5zkSm3peitcPOOVxMmSTyGQK/TD
AmDxlJpvi646ykkBJvTr9cc4gK1kEpn8YXiymsZuSsgWNk3cIPIegSdIIyFGATrwlpaUY3+UgWgK
fFonmfwcdmYcH5BDGS4q9VM52/6vhTnKPvYl6um/sH3wB7ocBUQGYCMj4+QG4/HGZlNVV2pAvlfY
OrhKFTIAgzZ+Rh2G6nzyLMyM4NXK93ffxcUbMiLG13rf/33qrYPz2zwVB0fzoBgR0hBBzpmOjC7d
ikQ6SWRu6Vape+naNeCLpsviLgX18tNv3WhS8RRRiydfjBYTFb9PmXqwYBKICWZdbM1ANVbAdiF+
jcc9R5txmwbjVK3yT10P1tMbU+TK7rCZwBHdg++HGeoz+RI2HdLvfKXYU/39cewqDH7KnwYxeHZN
IiNlSA2FgXWb2VIPzrbzRyYH6EdX38O5vXr0QKbFGxMV3RzKlPeuy5fUEOAFvi1No8YxeEzKzGbR
6IcLLpYcfk01dwrWtOC4p9HzHX5ZjMPrJdexwt5GurbyCcVkmTLH5Iz+3bvGY2/OyywKQodO9B5L
s0+DXjbbDt7UVruKbvVUDYcxr+55DlkR5w/RLMHHRbmMIX5cSdoZrP5mmBDysuVzs6fbOe/mqTjT
PKhzrZYcHXBeEbvBtH2srHV41z5353nvgo5ftnxxZaX0GqGrk+v4yaABPLR7LErzRx2ngzbtz3YE
mPYeSmsotQNWopbL72m4twF8NsY4mzQ62eO/5vjJRQbY4EdjRiAvTiqdrvDYvQoAMsgfoY8prjPv
dAaeZL/VkPZaEPQDlS5jHiFF2WRAqZHguwVsaTQkdCQbGUvZPTbyNCJF0tUkSCUPGraaWg4q6QPF
iB3Gtw7NI5bDR23wfImqwtHP6OoXzvHqZ/1PEnZyL2fJSKrQas1sCenmNwGdlckmgU0tp+nhCbmT
3u3Cki4TLYXOMbIaSPqAgL1yZ64mZQHw3tdvbEa2SYUaSJn4f2hIvT5ypSEmP6KoZu1IiUXcFIEb
2QDX/CZ7ECxgi2JTbjg3XZpCX+lMsAekkujPSFl7bHMyDTwWYYYiB3WadEgRanfnP7umiJt2xEuy
e7arDQ9QSrsRao9og0xpl0Fr29bvff+5cz82dj4TRJXuxzKxt/o4svlYxAX9zzyHbkGvtwYgpNc4
NfNh6LSogK8lTF7mxxE7xAV1/k1rxDTxCutUs04GVfx/dA2Zj6uxfidMhpDhKRxZYOotxkZPfpCA
WzE6s95qWJ/ta94y5w6+nfP3JmVPEkLu7J3AOukng0TW/uAKpBstdrVK7A55NSI9rtu+CQGTtYmc
/Gq8HcZIDUZxSAqLluo0A/FDrijJNToNbNnrF879ZzGMn1/DTCO6Ih9gJlaorDYF5Vc3QZr95ovI
9pMoXmtKjdMag0QSMB7S2SIEAYKE6cm/oujK7TwCYv+xNAIoKmUvIuD9+yjnKPIygbQ1MyLB6gkr
NKmxtMwVK1BF7B/nI2W+3HQPcFRiGxu3YbFodVkcsct3XVwt7dZzHKmA/rXPzhHuBlDJH2eb4S7R
W8uQnLOGPEbrLPnU2atJbxMnFDLSdTFMap/vVQbUBB/Taob6Fm8vuV3ygnvCMfPJ/bP7c2vEIq7Q
4LJdiSGK4wXa+9gsg020zkV3GTpuC9xJ/BtkeA5qNXr2uJ7hRzszM2+e1nSmU3c4oJZhMAuN7zVl
3YPOqPVUVWxIBTVJv1hdROGZ8wBZ/N31lrcm/sy64Vovm7cygYxugZD6dnPrR8WZk6e1ZiqkBPpF
CDuWEvieKW/HsZ881jZqjzWV+YVDJTJdU18gGexlh34aGvrTi/QmoUFklzPU6U3GGvtQm+Ed7AVW
ODnLvyQXesDXwhJYChqbwe9g4gdfv9wVxDzuzSliwnWcZDyVWBtUSuakQDqxrzQVBipHp5qn6Fmw
acH9Hhjo4r6mVYgKTZbH4Vqup0+hRnyiJsB37qxP6yqrm24V+30TnUvxxYZHh3wAZBL1ra7n30pK
bl91gwVzdWtUQindGmehhkrU+FB2UThA9H6qO8vadaLDFQXuXWoGV446NRmLYKeI2fKkkn3VEVxG
7iNepbQ85cyHyfCM3AAxN95WL16aRStrsJqd3OEdm2MjjZHGh7D2mvkT663AEjZge5vFrHshiK07
NIc5fBVgoN8EV9/pkRmvPRwv92GTAAvAlgDgYfqThHEt+ELNauSsfUNwWJj2gFbA5oeXJfzmhmh+
79rcYbYq6rSebYquWs/sOscsbPHfrbdEjk5M2lKVMyrURpJd6fily8k0TKywfTpj8j0nir45p90n
424BT42tLQAxaY/f946y7pIhYaLglPI0sD+dB9ZpORflI9xv3Zy84w8IBnDFyS3uPpyjy8AINH0O
UdmUR6QPqy/W0lVju3QR2GyDmqzqmMOtE6rNcsbjC7frHh7rYDkXHO7yAJDUXf0eFrDCi2OsGTCn
jZQtkj1DHnZXD/D6xttfziFmTp2MUL67tYg9QgO4GhQVtsaR5D/ZruLPoPBFq0hQL7E8aUic5CLQ
8Y5pWDqRIwCpkM4GCvfqf0zWYdmEyEivooOIeySEEAeklUSCWUSAqL+4Qttn7AEtTyYaVOl/OTkC
jh+LvdLmRaaQ0Gpf3ChgDsEUmEGdR9jl6OZM4bC8TbycRaMR8S0O2sebg1++RpsPCBaI4/9R1/Sd
X/tMqBeVjS/WceRPYU39ozwi1ke7omwXIHdVPTXAGju6bqZOqmWSgpJhG5KiZwAmeWRDH2Xf87FK
ppuMpOiYIgHZVowIEa84RVtnGTT8tY1J558/yw34YagAY50YI0aDWZAHrSkm14r5QtDAaTcw2L21
flr9FSZuIjD/SwZlOL1KONMrUb1W7dhnodOHaTaMgKNeJaDERXA1XfH9rDkJAHguyBpuJRSLsq06
mH21xMGyZ7/5LAkj7zqKJFfL1OavUf/fUqBOQz0FDY/4CnIzQPiqkXQWOtkAQKhOYhLwdp48GkLk
zhW/DMNqF+BiWhHO4gSVg15Nc4Nnl1402PzF70XiZqjWRutPpQ/lZcAAli2SQb2i4lZdM6z0vIeB
ipL3KK5cFDXufxV0LZWeXEaTz7vwcguCPzQ7zWNZ9rjmmgUEQuQ3Pktl3j+6KWvPeVNXySJiy+mP
j6pDJgYz0gFYGPwQW1msZZNV+Or5bbVU/BkhUDNLQ7Cihz2RYzODKc9jfiuQFOF2aQnONRI31PbE
9RT/NrRY04nylGx8n34iQR+O3AXFC4eFrqiG5ZgZTBlgmF3umhH++xP2qaSkclpmzmdGWWKKPyUa
gYfwEMmdRUrfmmxxRoGbkkQ45yYWQd6DDLuQf13Y0V0nWIAr6Nofsh2K+fnyJkazx42aeSWFXSSF
5ikR9aEUx4A+1rEHXBcoQy3v3P/gmEvbCDLDBtfiIyPP2MAKKOCaERwmYJEU811bHUhz8rzmlK18
xdyLFeF9p9gyNPKOcNrpXvOufS2l6M9C3qeSNrss2EytJAURRR78W8DXHOCH0CmdceUVaQhTUcrF
7AU2p5h46vC6Fn8VLnodg/pfgPmcTFLhXfoGR/aaoEWOcqlpHPNt/OHiwIBDsOe15ZMe+WQSBKLc
oIFq6NmvpJxd8an9z2xd4ajn5oU9I82nD2yefsgLcZvhrdIsg4M7sQpWZ0d3Ye/fpGByK1EOjv9+
41rVXweDsxpWQq64Wc8t+yraka5XsIdVI+2ZKP76Ahrh7kZJBhC4G675m9lHwxc43KM19Pm1rO/9
LmqCOa7muARwh0EEds9PdcqLTpyNNG9C7cSAegb+bC78xoxOrZoZt6dFzQvDz2AaZwe0xKjONNb0
HiSkMlRC268TC1gpzzHtIoFDbaEDl0ZYZjCBVWGgd5QNaCeCFDlwGCvQqy+cr879aS3Wd7VQjasx
iA3dPUOQItQB2wqc8oa+uWD0ufChg4e1R5M7MAelb9ph/4/MvG5da/kSaVFs0aKH0prkmZk7GLPH
r1e9vviobBGCjKieaTM+G5GPhxRV6pymCyu05NQrN7ay5zo+/wHkMDWVsImngjfhbtf1bNVnyCWi
g7T3cuWIuB7sjQ5+L73eDwYVSFi7DDMJsPt+qdSzbkdQtOrvtJhR546qF9d8Z6easa62FPpdkMqh
OLXSaUJHt8bwIguFPA0M/5iIC8MkGk/1wvMs1ni0HT1e8CEf5yoLj5vFzEPvVvNri8ZGwaNloZql
92CKqRSjjxEUM5LY7q2tM2WQE7K03LUncu50ssJbIpSgzGINKmx69+zE/uRHYL6/2C5K6spYsGye
xW1TkZRDeCc+4FtuO/kIZyLUEGTcEJsYYyb+lokdp7U2TL56Y37c6gEDTGXn6KN3Sma4+zABmmX/
b0ermCb7At1AtFXATBhTMJtH3ISvGx4qvU7DZol7t0jyUKjv3anbVQyz0449Bx1TEI0ipFuKNctZ
Xtx5/7Ml0hAOcLFfq83QkgpABmmiEdRadx979sHGnad1dXYfF1BuAmJssEusjXmdiex1w7s1MxND
E4C/6TfzhIhe0Kik9jTVSOf+1LFjcfc94LrYhQn/FYc8Y4U6VhhDxf7tMbZH26Pff1ikZoI0M11w
aOe6bFE43aiZ4eFzE+5rxouwwDGnXixr9r3nVL2vzfnGeCvvjComsvxKi8bPlwXXjmgyagS7gmYb
bPY4pgpyX915x4K21glGr24/ZaNy+cmpfukmWguJNMjZBRD4Nii1m7pCbjSr24pV2qzvOcd0AAGA
dWOTuWcvDgUt/Rt443Jw98NHyXDVv96EiZ7uLobITsHckW8xNENAG2kPayuSlRatkc14xEk9mik/
ctXksHDVkVHQ31z0fOVJouiM8sWPoLiJWOFpvjuaItQ2QQ28ooEKzO1cIjmoUmWJRGQ4IzAk9oEz
C5XkqA4QcXofqhdDOTuy2Ed+oCSzi9+ZDd1UQjvKSeSJAB3YU8lyyqXGVcxvGksEByQlV6Yv9NL5
WJyUdYvXwih7lV2F3L0M6QTwBNz7recvTQa5wD1Puz9hYeKAzkoMy08xQ90/Bh1LPCyUG9UrvWaT
/dzXpB2f7JCJtB0sYbeMi/EB/wtaJ2jJrTY0MBKP/4l+i45oz1CI1XTRmARnBFsVlsx4+SAIpZIl
JPWryl9gLMXoAuZPGXBcqZqq7s1wjg2MriV1ooE83PV4MbTfK6rRddXm5zjzj9uu1wtxjn7nQ2Bx
gE6YYu1Cpm0nR6sMWHivAfGmrfs0fJniSku64221EhenxkwFbgkyva7g70ayNJBCL7a/syGIOW4r
5lsd+qVnaYIFhgpdJ4yuavP8NJJx++Wvzn42d8q8PpTNIJ6XiIaS6koA6QYs69/iTdZnX6hAUXGM
nkw3ezLJ1XFPPWb021soI5pmCoPSCjO74N0fNgZw4I2WNvX39msQYkRCJA3huVLxJjLb8im1VA3p
GemOYmES2HnHKZbQUPg5mQRIWr5DkhjGwBDXhicwEQFM4l0o3p9p7WJfaJIzsIVdTQ+HJP3L3ybC
jFGSE9ABcf5ux7hbYU2F09EjPxZUaBexM3IXk9J057FTZa3bwD9Quwzy2b0F6FegGaC+L01iLarx
PXpmcoIYC55FHfHQPfcT23rsJ+QZF9CYoXD2axdmrR9aKIJrjHez/veELNmfZAO/emP0In8a9FbQ
bvOlhJbQKc4MucxWQ/MCZ28DWQHdJn+qO33rfpm4z3rTVFJSwwUpOg80MDULSm53pKmBXYeEo9cr
NG4NkuviCer+9n6DihwOwdIYk0xrU3u0O0vIsf3J4EPXthF0BDtoikalnQwOYB8pIjji8HS+rY4z
FUXd6GxvN1MJvra12ohC4b6CHvoupJhd5VCiO1OAkJMYkHTWzrHCEcUXNACOv6ZSmkqiODrAep4e
d9WVqfUe/58WUIWUxUNrc3S9/Nh57m0CyNgSmuj3cl8aEMgCKf9P1XBvpVQfHAZHr7d0iurhotVF
50exALsuRorXEgvsjHE+Ivk54eY3wl0vyn9fummNwBwEkyQASbz/VE/ARtpzSVkJITLjTyhLWZBx
rWHU0Hk98LZufDl3AUQqfe7qL6/CaXaQ/3Fh8QidKJPbyiOUjInl8+oH76rJbmG2RN+7PixXW0RY
2BGWCoTmYGkgaEF9rnY3a9hM36SGnRqFEoRwRZByjOdgfySYfwyGQHnwYfX2TjwE6u9wbCxAfMmx
W+WAuj9AdBJpRC6l78UN+fa2OEZnRzyjBKEIFoEVaiphlOTCJrqMJIWIMQOkYA0MRBpdF1mEXL1a
qzeOpRa4Y6NroJgwqt+H/1NwsAwDRbS5QyVo6WPkQ3ek/g0claDRy8aQ0p2zFvSBN38nQIMKGsTy
h6eGWC+M8itewoO2lK5URlBWhh/IhzV519YCLxiYE1iylwHMDdl688GQWpZz6GafMnXFb4TQaW1o
KlmqoCCujCOp+XMxuYG6fFdp9RlrymW6UOuka7H4luUPKWriCYJcZ1bpFicYXBgK3nOwe6idd0g2
M0U8ZVuKaje7ygK81+Z/RJhOQQynrap6LnKzlg5z9K2CJOz7oouoigdi4c0TBdOxrTfjwettmqrj
X3A/qVzu4LMvQp+H3dZCHIzJpsDZaca1HHdq5mlE7kIVm5jnUXgWKQTjqMQ4KHHeFZ13kADDUzVG
r6S362V3BM3BSpDR37A73rgvY1Ta/KiozCyt7rho/7XqdrG0XZ7m0RK3Wnh0Ga7Piq1RWzmzUiij
aSn68FKCKUzvtAybEm8BKtsNu4FJJRGeksbbaqSuyRyrDx7CkEFPKtsSetFkLR9xnVR+IQdXXHjO
Ty4yRx3MV8MzZtaRLYPP8uGolqOoN3Tk5frjhJgCpXl22xMXNf5xxs+jMG2724hHnY+jXlb4W3th
vBbkiAOH94Y2f2is0LZqB9C3RVnWq11FzFMri0LvHz+ASa713FbTwu163fO2HRatE2X2/6CPHxID
PSXLyh27QY/fNPaJadlN9yqBeFOiiYZWU0FCjXAY/83loOsvXTsUJlz7cRswmOpQNFp4/BkIGODz
RHNJYW5/0Lsmg7015/lPtVafgc73kv8UffZoPldnCUpehIDQ5++h2QqDhIobJh81pcyUzJ+T1o4i
2q5+Jxica5iqSXFFCWbFUbjMCcZ/uWgqcCg/pL5d3j42Kx14dQLDaZ01AWH25jqelrwo2IDAu5cp
ZQih0EibtqajUnxrxTw2M7urtMIejgN633mvYLwIoyR9tq555cS5WI3EpKqWe1uAUROMgAoVEz2X
vjAXCKR0Un4Ei0p9QIJKkcZRTLzDCmWEfzgu9UjiAVD+1lrufQrh/pRVfQIwKVZfSYgTVxoD2UN+
Pu8zb0VYwnYyy0O8FziFSZ6DOdW8Ctt5z6VLvZrYWLiK6Xj9c1Kmo6rYSQsn1IsFIJEJ89Rm3g24
Zj94thVd1QbECgazb0IdklHB5VvVZNEhAKYROKgZUUFLnpw0z19NrUOujrmg50K8oUoQGt652hkb
aJxUSKyCTFRiuNTS6qsh/JAB3e3wJXW9giHDkynx6C0cdBKcDntszhsQanmA9a2QPQ4dldp3/eV/
+qoJEsjkXiNsoJa7/HoTVe8iEl4KuhhZd70GrEzdSsVyQqG7BI5pALqprEM1vDb4CH0xkb9y6+Ux
lIwD/GbURVrRDBRlXidLt93euSBdYWsfnjyNUhOVvBIA+yt2iDcp0TgvCLAkh980JR5qgzskS414
EBMTuqBLIagPKG8LEF73ASdCgd1tPyHKL22m8tkMmAJMDm20d9q46Z1bzdNGJT43agxEcubFUW6S
FlwAJzOlfCf2+xb97/yyFXlfrN4qkNg5Z8FUkvB6GA+Y8R0SnwgdaUUc/xFyGSNJYE706tUFgdH7
RM5doZyX4TdtZJoxNys8cDXogW7bkEk2UvdK7nIxbHBqbScVdypnGGoe+L8vKNoXs+ynIQLiUdwr
QNa1KFNKGDlA4Fylf7ePLXmOEb/uAsghsy2hW+Z20LSMrqgde5aqfZQP9oLvdBbJW0jZdwAd7Z0+
KWHeHDyzTjRh17t15aN3P/cvHcagiV9WZh1pqtzZHsIGMX6YENVrlfvIZbB/MfV9KY1C3h0fQNdc
EYchiyikn+f42CDILCuicvOQr3yeBGUkEUrIoKPzYL6/5WAMZrQakjaSmE5k/hrC0+RVd1MHPjui
s1DmgPNz4kbY/3dOfsSzKSKITuH47bhvfErv3fD9LwIpb2smo6gU/RIqk4W6L0FTb8eQrs8vW7eU
fLbgKeTqoq8y+ewFnubho9+LwvZjnDQ3PvbTfho+CkGPDlF+WRhn3TYox7UeGlh5Nyiq9KuiS3nI
e3XkeoekpS+5tnXhJh735UppcoUR2JI0PLeuFO1jkvV4A7VpWu+9YvPemNj2V3yGdqdWkW4c7EiQ
bldh+eXtHpOELizAse6W1bR068dkw05UKoefj/hvpIyGLGinqPJJJwpjsbM+IJe51VQBBJNLgSFz
xEOq00QglNrhh8Qiiiod964bvO87mQfp7sZ7GPnZYlWrU6U5rkbdW9gStUE62lbBZ0ZdfpHqaiHz
Xdb0GJZYf058OsUYSBzUhoiRGWZHoc5Sxnu95HSSG0f1sQ3IEwrtRnRUUg5+AtJJiBc7P+xCio8C
mF7iPonnruDZPFvOxedChtTjBfqjigdR631dP023MKfsktWQh764nutYq+BH/WrVsMiI4HP0MFqK
KeAHhhXEsud69e9UEoZMWeAtlIm5WGbttbNV/CdBvHkK+7+brfX2xqbZHjiwlGerXAR5pVkkGKO1
LYa5omMQoanzIJqxQjbZANWAzNRZ7zgBWN7nJwSeVD0O24h6MHDkzDd0h8hKbklROLw+bobjDYmd
uSaD0Lbeogk+n+JX84vWoUjJv5zqAR4IeKboUaEDKdQWNpa7NNheNk9UhV2gbcKwGYqhvxZahov0
kf6xhOJ1ybKfiMwzR97niCvpn6fqL9OBRsGOpmlqBIPE9rPpn1G0I9dtBjO7DABBcXAdp2A/iE1a
1B9Si91ozEVdcaGiseWbAfwGk4GBIqf+hnuOTKcg4rr1toyNxlVXNRnPeFZmLRCFBitD3eAbmYYF
7HDud/oAdMnSK7/wk7PI6xQD7y3L1RELCk4y6aTcBB7vkyonBrIg54XoPeGgSfUjkqJDCw0lU93g
I78tqMnr63gnMTcl1B9YrmZ93pQRolviVOWtX+AOeNvLlp9wnreq6zupvRhz/9JKWBacvhAIi+6k
l2BBGkaiJpGuP3xpK1RyzDA6a67JSFN9O4qfC5a8gkOg8DQSXAkfMPwBD4Fnt9V9j/oTEuPr5JQ2
i8ecW4nC2uXBwmUeaSKPbK9VQ7AWaLvrHQjsPkRvsaqFGmKyae+3b9StuS/OVF4YfkPRqNIKFOhc
IXCxUcsSwuxAZfZt/lq8ex6oqDJH7esmVk/STKoDLpU3d3pv+HFzed5kHZj65pvW78VHjnQ/vmsT
wJtFbK9CoAuC9TVN4u3WyTxOUVJBeZSsIZEoIKmj3BhVcRUCI9uUy1HTYKe/BfWdiOxFAQ+NWq57
G49PdUHXKP5iMTpi3BwHpiK4aJ8cFymblu9qRxUiyV8z5zD1fJsP32yOOA5/EvGomcWhqsFDlROc
pywnXPiuasScfaQA1V0hnYgb+BBG/T+EW8tyw4tCLT8LfkLxBXMDESF93VfbHt19PZklSeFfFiZH
oEXyPJ40mzHCQdC/5s4aZU2wyTcDFcpXr52CCJCEbtT9dVVWFy+pWskePO8kBVKfsg6RaBbopowM
p/GOsHRLew+fO+sjG97AX/SoI24XhqwhT8VE8P3Tn06qKCWkASrXe7p91xqsgUEeqUZvdqJVBFqe
iM4h19KIy3Ud32ukCxXTtpNQN8wm5++bh8l4NsjtGte6dIaNyhLG0w55GLc8CAD8SZZcEFx6eyr/
yfXnnupN6tHW11VIPy7D5Epn+yqQmXJeIEuLoCQt/DDI9Y5+0ON4t9LB8vDCLpO3DLOnAZWJlAiV
KcI3OzwPV9nGwkq086PhOzumB82t+vGSh7C+H6Cs4x6070lCS5pa5xMO8LPs/naNFbumcvBvG53o
d8NegqdiP7jxpAzRIQA2h2AKRBn6K5kQTZyaR/S3hFq9PqAIHrcitKoBWtAjxQWzr0CFbDFUyW8w
FfUKKjh6VgKfN8Zr8dXD13jSxZualo6yhrubXiRAX7+Mmt2SYnW7JquuAXiCjqVLYRrJRXqFZfsj
by1EopQCmQHaZmAbJogFvhJQqp8xfjmbnesZpCklnbovEmYFoOeUivQ5vMbIWmRsMzV674Y6IU3W
SfEeoXf44frwZhGOsxK3IVukMxN6D3nGoAvrSM5O/FKIuUPxMubpeAZkSWNQ5xEGvNLhmAKngXCN
2O+KKYVeaw+kUp7LM3EhxfZbqBiG6yyp6BfNN3rI1QloNd/Ng22bHOK/RYZdJ1tAgFL3VtcJ1brV
ZeMNjIK2gldpFRcNkdjffnz/ndnGbD02lkN0g6W1vCt5nAE28AR2AiqxoPNgj9WRALmmFXSVrjNz
eQwk6Qvx5K/bdM6Fh7rI3XtVVWpJaRQpAFk+1V1BOHkdvU0dhJ6yx6Acd4eoOsgSARcXT9tqx5Sl
qebyyNlMjPwHlESjGxIrJxD9nFo7CaTUHtZU7mDDcyTr/MoDXBZyk+kpRg8qR3z7PeO/uo2b4s9V
DTjc39gilsW7s+Rm3CWH4dAcTauICO0Pq9dcsgvywmNplWQ/6h33ZveI64Sp7yBNpoDjOzGPVcra
l1DWvXgfk/g+jHLH67xtosfInYNh2eCZNBxi7XYtH4wS/kv7QRCnsuZ5wRtSp2J6Cxub/yt9kmdf
i/s5xljPoN1Gf74q2fWLbcZWMXwQt8l2VbX9hR0MBvP6HhIXpYGRvtY2YC0cPQSvoge8iUC94/Wx
8Mr3WxAztV7DDG05DlXGbEaCg26j7BP50wHqix+1nuI3TbQP2DgLOV2qGZPzcD+TM1jSRcjDiqGX
3WturlNccKofhi1vH7Whe8CrmwLeiO7u8XgaWXAn0o5JmleHxlwYhwI0l5EJTGVZ4crcXDcC+PoM
iFUCooB1GHdTl17izisZ/9hnKcHyzVdd3KQLImA+VpSmps+X0xhBykC5ukHifkx+xEJcUs4i6Usw
ngF7AsXLyczU9l1naYtJASgCO7UIx4xtbkXg7/cKobw+CrOgn+CT2m6oOD2ImxifZiQFqLOnVr7a
nf+BoiwhJI6aWjFSGpoXg9fQpN8Q4Cl8Xb8jL6PVTzodfF1SVTsd4CrO0axC08MKd4stPH9acaAr
ZM4gAu4RwGH76QsiB8Ra7SuZ2PWcZvgfkBzDnB9pgLOd87sJWVUCueoFFODjWtfMYkynCWd8RWUX
z0nMMJirwD59wVgy42AU30xwPE/8Z36XJDonOTkMojEUDRHqk1f+Y0bqc7hwonh0DIuLY8u+mqvY
wEuK0gUjhNR9i9fy2F+Os7sfnR/cN+PVRNOIgmAN3kuEaEjpw0AtbINXdhqyTaknx4Q5KeVKH9Q1
e7NTbaULGjU+BBhzLleac/VXauumD/iddLdow2tL0bTO+uvODs6uWK+zVs6kcJm0fqQinIdKq2Yx
NWk967XXyYkyTy4Z2h/El7hPImVu1cAHm60SQ/x9rtIcmmQkeKnuy5cuvHZR7nXirE79xPiKgWi9
rAzbAHCDm2VztJ0H322SEUvvAdIAsXPXN1MIClTjjLCVB1RAs+A57lv7l4AXHiAsRdlGhcUMU1wh
8Sdmkb+cS4CiOQ0Dq8u5iN3Oi6lVW0Iken+m7zX/oShbCmvnG/YQLdoUVKQPW6uIhDyLVv3DGYxL
5Qzch/fJ9OymQA5U/YAJRtO5CsHVvNxEGL0tMhhLGBvMDa1WqjzN1Zra2bJAnoT7QtrQxrU6h6lL
32hMjE0ZbcMwGZQ5hxJER8mtJ3PrudrGbGVk+Lijpzmd3+jq8NxojFmrZZ/8jUKxf3Pl0Ko8Jrid
RMKyNrRVogzFLEz6QrcdPWMAEckhHhqt73MGpaep7dsfpfD8YPJjbwnFIKW0Oa/iVSfY8jtkBPfH
d1ZbUr9Ph3fghMDTQ9WRNFdNBGLD0HC+zUBIQ53UrUCh32stR1AeN9a72U9Eac7NHHY1RFWHi/Cv
lHCnqJQIo9XWJl7LfXTov/xrpg7odDnJc1uqfgSvBnxVd3UqVeZOM/ujVAz6kXN+fruoIuz+6GIR
8HpcMy7DQQV8eg71/f/FONmUr3yqXxmoL582Pbg/tnrFOlvJbO1X0+8pCGCHmDfXiKUqVRrRcihx
f5nUiTo1WE0UQH//I7117iFfLFz1YmSPR0+ydXk8Q77PYA6BfoW5pF7C+TPcbbK8rI4kVZgt0Zvg
i2Q0VD2LwgQsHLdiGCw3RjM3ZfJLX93OekImcT4+l4QK7qhWws3i6aIyTa7OUg+8oJ4D1D0PUhC6
5pRyUNRkGNsNIOB0KoVHAx90sm2Q40/n2uVZiFv7clrZflhD3BXgZpz8/0bspqQScqWgh4yEYvGB
XmK2WJQeRqzvSuFRBf1YPWoHcr5c07n0z6FrADb5DkTy6Rxp3FsKR5qFkCOt6sVKI7cIeAjOhORb
tik6HsXImf6c6pui8nTqq8nTBYCHRO3KO31vmIvmLKwm5zMIVrRkKKuG/UQm1Mz/bAmsn8hBpGJz
Q9NVyVSxU9TgXu9nA5mHyVRVLgqVki8kuJF89aD3vubfyy03jz3FCacMRVr0yRFvxvWzptXyAtPN
WibOTNDMofL7xiEDh9RjshwbiQlQix3CvLzBtaYWXvqe/BM6eOPdKOD5wBfxE9bmuOxEp1WMahKE
zIrB2hCSUYZwL34ncgvMiQgMULg+qhaQ93M05SYZEMzO87NIGleffSz1PT/McvoFuJWJkNRPbU6o
FZfVD4WM+J3Zu08pfk43vgWrVsukzEsKnAmdg4JDXZCVSk7X/0H8hBT0sFxFNaT8xVb2FwKkUTUX
JluquUwr8TPt6O9KehFScN5R2le/RzzHYADTFHX91OuYT759td9hSa1WyWFuQIajHwP4x7fbLN9p
P386/yG1IFonWRUG9YDU3rKxJ8TValWGHNDszI98alIV/q7MU06tLEzPLAMZSonRDbrONEGPxN+9
Ds57bN1YCG4MOnotNFJg+CvTSZd5UH5VKn7v2CB11H5/FuHdp8GV9q/xFwcrH7EmFv9B5XoNH9mU
MOgFeTafeAwwuEmQd7+YvkNxWQ9brECMSXtqN2PQkxmoM82Pn1wJVnMJ8SF8yk/svZsalh+VviAj
QZUm2/ivgIA+k1yYgs0BhjnQORWzmiEaQk6/qDl49vJ0+FIuJR2smPPRUbAIoMroJZR8G9KkBNrz
btwtiepDVmRQb1o7t8KICtetXAM5byzbbGwOJaOUPL2SgnVTITCczqPQIrahqgnvbhAUYquYXVlP
uU68AMJYMWXfxSAIYuHci3Rkn+eqtVNFyydzIvb4qGGMCcfBWjUyey/6a8UFGhRdu/KXKW11HkvE
mFibfFjTJpy2tw8QoGk6ffRpdslXAZxCn7/bs5ACruFVPebey/j78qrM74orbhTThxCSvHcDiThH
idLSvfywC1zEJl7DaPLvT0Ok2hr/wulGmPUE2nFt/0RRjFng4CbSatw3H0HoYtaJSfDDm+41a0oZ
0bWoVbLco5hHjxiIqpfH/MYe5IwvTtS95HkPbw5FKR6V08v/hgB5I2AjkhbsQR95Wbc/Cjvr/fVa
1NPU2ck+Op4zXhCQnKTxnZ28vdzP2md02x+mfe1LjHH96zgByxBF7/Na0Joc1MtXDcKBSpHnTS9B
keAPUzy+wMNXW5HgsmVYS4dFDnIawkxBTJ+pcwPZhgsaTt6jZHMtcALNgNtDnbYIJl9Yk9pdXG+D
V+79YuDBUmnRkbzzt+A+jag99BBWLqPIE977tKBO9K8UJrqLWi0dhrpuzuDAQ1yS69nFbXd0aIa0
dFUO9rhkD1DELO/P4UzaBFb5QZJenvrxCBrqypNo3dZ3XJ4Y0XPb0iWtelqUkTFgrlFugN9M12pi
pv0Cvqe/tnfeIH+TDi+6pJ7FYJaJNUEsZ0+GQRXifSA5K+JflxN5yW9EQQg6L7c/fDEgyqf59Ecv
510fgRVXB0atQW1SVRwEbqkfUirNRw5e725emHTTg5Vl2gQqGoddLKlG3wEhuAMsyiX2Litd7nY+
ixc3UW6yYkQMvRKjUUTIkNBkjIjvnS/1eQu6cOM3JmbP6a2+urj8EPhu9KnWd/oSL6zMEDQ2XXuz
hY8QQmGXOAGB3VLz4dlBITQo5jqGkUKYl3Q5sFSN8fyCh2rv/rGtBLkaz6uco5V8jdYjxGEcMU8M
otA55mCrznVTcB01a6ME/eZ5h0MYqIfcYTGEYLlQtJF7hTEhwyGCu+j3fg+EOXlJN06fjaoYwFfX
ahx2MgTMcdUgb57J9JK5ehnjr5sJvLPXPyjyC2CUEPEzMxb4LJjCwwLwttwVU6SPBTuQecAgOI1J
H0oRSqfmdNHUrO51Z01rlcU0bpW0srrS5lgRkKre60jQT4P8K8wRMlS0Tcc/IIUdX1gKsyfXfNO2
YEDOL4zrTdkyAuj4Dlzg8uH9OKLWm0YQjj/6DAI3XYmxiiTmvirzLEJtxtTDDx0SW1Z8TThW29nL
Zakea+BKq4LvckqcJSwOXsYRUrEt3TdVAbl11OxDYoeb3VKVyAYcbSX7yVgFthB77oKRTvYfn/jZ
VEh+fLLPaJQv/sxaEPq7d1ST9AfbtBzvW3yiQIi5MP7XNlcSTVOeC2L0zwLtgvZGK+Dh2Xv+AqKn
BO2jqjdPnEG1e4JXhF7DBmErVYI8ITvbCYlBktkKsDsHZ0EBcqunfENuyzEh7WkO7/RMqVntrLDD
mgrtz4l/MSe272TF8NMDnmjRw96Ht2Bbicc59jMEwbiUmTZZymSgNgSEJNLBdCNR2Wi+5EzyFyGs
LVPa2mFnWV5+ndlnVTZO44Ldiiefz4j4mJdGX3S0R4mJ/le1U46VOruB8UpXKkQwbCCka3T/sbsh
/lTVs3MYTd2r0mKwxWD2FI7FlqXBBk/iKjnxzWp6v2epSNSR938rXW2txRP13OpLyvlOdVZMQz7M
R2Mi1C00EfiUo2y/a9tNXxyqHOvBXan3OWEppzmo8Cx6qGnzl9lXHQnX8Mtd9H429N++2GDoA1Pf
t7H2/a/dR5Yxt9i4JU/5Onu2CAccrG892qTAH7YNQeDJONtlk64ZygOG0rx85OJEKMIrbBAy7ppJ
yA0VcP4SNOjw9frSc7/LAES34OU9Y3lTOhn8Cz+sH163wo4/O3Lw1GXeSTSeBO0IxygqUnSS1pZZ
3cgvtm0qrqmt9jux+RPV7O7bMknXcr/TuSkIscqDrCZrGduZMFlfvbxsOPSTq5UkiVfOOmqhMNED
2YbKLhdIgN2gaC3lcQUuKuHUFqfebAS9y3OzJUYM8nLbuIcyAj1yNarJOO7AEDrYxumiOty8m/E4
NNdUvvaZh2OYW0jOi2Y7bM8YdCyCNb4pQWBZ9e6uUQVYt4ZhBXOeZhPFkYOYY/ErpnXmCy4tpFl0
VQrtq3lZIoKh/J3BfUunt/p2g/Am+pbJO5MtZL3o9gW1s9+1eHX7nzc8syzU1IcrRv5K4xtB6fpR
mLtTTn9KifvTCHaArtlK8P84NSkYCuO26dIrAZ72mXHhRrDDpAGc7tNyTqSMlHfyjf35EMT2MxMt
BLpHZTp5cCsL0eTw+X6ErPuGDOMTiJ01AYHsHsOECXNuC2oqf03gwvrKvbJlfLvrH/bBLqziDMj9
3lQ+qYhfoQL+/h1LDmJ8E4Nid3cJcxt3qvRCpyboPpAzs/zhq6t3q2QHkuHpefoeGzXDas7r/hn3
CevdDQPknLVLDDc8obIV93lQvEzuCbgfa358jQ3+BUiB0oQtkmkSkxW5ZhdHYThZCeB7uSvydjIZ
zCBkdIZGBtT2BN6hnfCbmbl62XmSQ9q1uYWn7kNi+VEqf2I8Y/azTiE1p+4ivWFwaDFdMCQFpCT/
vJhPdZ1c0Ct7SEZY6aNuLCmDUpjUnWX7SOc2ew00jXF+++9E+Xu8jLV7BLQq08SbwZuoyQ2J1iSQ
C575m9sJKVwt2xolL6qOrnU33KsjQazGHml8mjQ3tuvNg8ewq+mEgPDppYEAyhT6g575xWHh232i
ZlVZnijKARJdVbce8IYOasyj4+rPrSv6GoCKZ+3TpUmcLNjCNwh8HPgWupHoD0KHttPkfOlAjbJK
67JfjE4qtgtQuiibvpKg86Ctd/MTgJ2LzbXtKfE3oG0j84JJ7j7Sf57sy5RfA0cmYoP1s471oMNn
IV5o+dtkPansqO6kIxhNm015jp6JG0d2+UE1jaQ5A3/bWqxRe6Pfd7LaYCGjQeW5blyThoAmCT7w
CYMw++lp2Kzv3X7kZ2Y1al2K5aVdM9XqaHhj3mROX+btSX4oJlFW6lJoY4mapbb88uohqqrDtAGM
jsPvsQHhwymfKx6U5ytyYPpfz6AB4iYzMDpSj93c0Q5YiTG+e5taHDbxJx/FJ32LJ8YSkqri9Dv4
RC8ZU1BPOCytbb6MUIgH8WCRLTBCHOZVO2yHcAdppVxFkxfvSAlZXulIH/8ZdVEWgS86/vZzaV/L
KAAXiOq1xdELGMwkxIx6VwrYJQHeWEvEq9CYZmA/c+Nv6Kr6aeV0glNdjyR+pxdMvAzrXr34z0YE
2Gtka3qluOto+AwbGOt8O3GWg7TxxNeUChv01LFBWgK8oWRbXG1MAwsxQl4kO0NfAshdbd+kWknT
FUWUMy4+Xa4cL/IKl3z8GOKPJg5cfDv8YW2wuPBN7vYRqSPaoc4QhQkTQJhbw16GJVV/Uj2JoXmS
zB1k/AMq3yM3Wlu3l8HfJ+BSmM3vOawWs7yvSIEX/6X3L7vEPqfZgUmJ6Cdc6g04NRrfHuNy6PNu
dRy31i+eJBdODPY3Unt6dlTGhISBghTwQbdQI7G6qy7yV2yQXGAZf6w63K9qBI+MaL8VdBz0tmMX
eEYOPFw7AypinANH2EvPVxFbUC9ERWNepiCT713VrbvB6Del1GbUVsQ/7nFsTV7FwLYeZ1xo7iF5
ZBu8jjB5WomzrTWYjJO8n/IFCliyBXz/tRF/yicVyuaTDVH/8CKTRXiUIUPdv+CsMNOJIyTpArs1
Kms/IT9WmOhd+LwPwqst7wEviD/+xTRu8yG9Z959WnumVIyBUWmDnb1NETjnXvDTimOnA4/gfies
Q19xcelmw6OkuOyWGZz9Dm5xEKBzbylWGmgP32UELfyzoJaTV21E0T4knpy6qb2l78aOK42iGvkZ
JeXgKfTCpeVo+5Y+Tqd7IcBZSD/xbcZq/7YiWUsMLys20CgZW4WnTDrYCWyVymzsFiF/oCs3bvWX
CsQ1VZg3k3AdyfXDSOamPPCO0Nw0pvX/RIbeg3DgaNFn1bVLLpCV+NSXSB0b2ihXOZUjZNQA/sqN
ijm4yovBChilB/ns10bpSGHEkuDgPWuZKIfVy00DGcevNtK3lJaFuMUvMJpIUgyXnRVngNvsLwbX
kpVmPGU8/koJRXI0IBqvfhjq4nUzVIvglxk+iqwQuEFyXidq/IQ7qlfL1qSzxiSOkKdLSM2R4xPN
CcX/1uRHM/O2TsdK1HzAoDHgR4UP2b4dn+CfASs9W8iRkwLC75OnMQCUc0E0T3qRHoq7DbQBZuTq
r7m0Zn3C7hWfZ51Rarxs70YOVXeJhK9FdiEfzdF8XMZ6AFCjkXyIIBTkUHozx3gxrP9S5cLg3COF
hB/zgeRqk/N6YtjGsaDnwPElo6fICDjl3LK3VjmZ0bVdkW3wCEMnIar3KpNjzMUGpcGfdwx9NeE/
cEoSMD9azFdnXcpT1WwcvHt2sqpqW3IdCctwGMYGI49np/+5NDO59Jpfs+Io4GHDEPyGNOhvo93t
T/CPJfcIuDVQmW0kCK/yyRGjXyKh1W3jMmz3O21gf8Kn3Nm+Ck5Ai9YE7BGKPmeKtgIcCxFo2a0h
DD0MsW8SzTVwNhG+djI18BabdvqJiSZJy814809ZHC7sF+8M8L/xs7xVVtkX0apNnWEVFaiUbX7C
+yVeCW13OzN1mxBrnHlNRfDjao3J4oHJWqCKx3EQ5fC2q8mFhU0lrHvHivJRUN8hDRGQE3Yp9K+2
9gd2SNNFYnoaX56Y02G1rYG4FUWNNHB1c5zPNgXU9Gk+R0VzZNQxbJ/Tr1khI9RdE0yZCbnEli2F
gIj5oMTrglWvkAqbuFDWTpIRbqWtWnq+p2FoeF4siRHb7csZHOg1ZiXs650X4XnwoGRqW3zMeQq9
D5cZCbbz6mB7fUt9CWbAtU18rmABG8sjac9On3M9M6fWb3MaQ/EIFIV+xvXXOh3XAVxkCJItdS7k
isXRTsfb+amYF2VD+58SjaExRVsvBlyndCt8xDih5O13wls/ZEAfWSZGuTZSLrFs7sCiMXvZYKpa
WcmGjUXgJ2uWdgqCV50oJL1ybtboEDcblRhZhUFYQ+7KvHJvb9Zls4w0xmTxm9OCvXkkIEWk3WsA
UVlLssZ23eK90Tdl2FA5mT9nJYT5qIBLu/IwgdtTkrHf2LU4ZqHbMUhzfscv28lL2AOhNd30GBkA
s6m62OyOtKQ0Z0vBRa71ruN0rHiMDGQJdKDtCXW8dvw61wyP5dqWNphwf/Fj6qitY6SV822rzCbQ
N0WzM1hP2CcUt6s0gm7XFnYCfRV7Ev4w6jqa9lKjQWIJAZFbufndTdcejBB5LhjnUiX4PEfCX5h+
VA3joJUU9Tsl//SZG8Lzu8XNth8mwK5s/0Vkhh0QIJRCO2yZLwFMbOOjZBULQzuwCF9V62KtCmRG
nGns99HMrK4JUTXXevW5uWOHYmhvIK+yJVvsTuUfQg7B7h/8zHpkELf2GnERWUMiBZFV3HdAmuWA
COqB6jb4zQjrJ/y+/PZYa6sY49GFaRP4AwEm2heg0WPWjg+xtITvgG9OQ5/ZYeJbscuBq1zbEXCh
IZB/yJ3sDG0EtLHiIUkkapn8wy4guREDmuEdzoq2TV/yC+ThJD5UBvwAMpKPBXEpBL3e/x/f6FkM
6sI548eos47JPqm1QEnquJ3YCUR3KJv5jcPpfjlxTkWIHc2dU/yPWDxZDxucbjLJ29MNlxZwQEHD
6x8Mp/sEOano8GRINBqCqmGyGZrWmKIZJHn1D97ODAbjwohoqGQInZvOhCHJ/jatVU9Lnqn4gP8v
FdoB87Xez5AUBnyijJQwETUU86xsAWD6KtQtQOqk5nNJ/78QY9PMzH4rZt5jyyzrT9LRZPpIV7/A
tb74SeZ91/KzVdqFypVuiA4vtsT7rJGHRJgSERCekXe24NUf38AdP1lM9zM+W8YyNPdKkgFhCZEY
s/2oYFmeTeanqCIMzSUCbwUwEMLyT2dRPFqfaUI3/40JBSpDju4ke+sjORZszTN9qh3mfBlGFsYa
3Nblnw4ycdisN8lsUoYS5RanY1ZkmjM6EZQvdJnlTmbMRbbluMijsUIl6/SWEgHF2Am9pisyrFD0
rjxu5r+T5TAe9ZD5q+tvpK/rrEvw4nr5YWm1qVOkILykbU1LMhMXrOS2tMxnJA5h6t5LPcmaZXQx
kAZXpbfpd+JcGXr9Qg8gnM6gcg/Hbe67bZFJ5Sjdp3n9Lv+l5Dt4AiQ5vh95MuZuu/wqbGA3EIxm
H/1LE3iK2H16ag4CmPNIfs8jlz8XmhQd7zT3QdnKxzmnzhfza2IBZSqVSWKtd/6h4H02NeOnGjKq
VS0ypXf5rcu7JGoN0+PsAvFz7Ik/rP2+2CKg2jLaHKTX1/Ex6jU3GCHhJBYsuYivbS+Jsrmfm1GX
N1OFYe1Zv0eRxh/HqjY9dMUegiOS3Q+weOFJvnzzKvLDStUqb7yHQvWlX+5H1XcPVv7/NvnqcgS8
/lCkB+2esd85djKXqlaO4JTuAsEe3PajbqYaoxSpTJJX0+toMxsVQIB6+PdT6f9jIH78bqD2cd7f
NXprQeeFkte9UGzFgDrRXolvB6nBiu+vTKb09fhfY2W9X/I/nztUEZmJiSfTalNWKZg/1d0WoXe4
E8dIX4/kSDsf2Feevc3yvxtQNhOXZKv/o2myNIAUXyPFxIn9FdSFOMu9iXWD/oxDfXGEM992u7m+
AZ8nO3B35vzYhRNA/UFHQAGjcdP7zw0mv6cUcYe68f6NIB/a2jsBv7cAEFD2BSZBQfl1DYUDDsvI
XEKIzXj/K8QLowuXgs5tiKZmxXXpbmcPlRf/GCbiQOs7avbQi9qips24G2cb908TsjPpcKYEfKgZ
A2Y6MobkBwpo1rhMJcl+CwON3rW38c9fKucePGzl7ciLppa/Yd95IrbnbtoTLelx1YlvAHZMGSeF
IC/x3riJFqYXUyt7Sl2V/mKTanB8gdlm55uTaAgFsVRxRvvCOZKaqfAPs3MJRlEd0GrsgNFGEuNA
Vmea2qxts+c3w1S95EVs1WKEXEYGtlp03mGxXSp9xMlb+6DG7MPoSBqi9RH1BVldXyMIcDAw3X9Z
e2iKg7fwEDrEUJunjtVzTJu54SB0atELpeKyf1/b4m2hjN6pFwho6a/XnDepwB1Gp/ZKxESWAI0x
GWyi2IWxkKf8iCUG0/rG1FDlCv4aRELe7dkfVe1Q9ctcpGaVNnhOe+J2ZOBOlmHwdwYYTjFAAs3M
+LOuD0S1QdxN6MooYvLEEDYXBKAMBL/WU++2S8hmae2NN1lrRrrTImcvTig8UBotSun6Z9S5Jd6o
DN2sWTWyIOtHzTOnZux0sXdHI//5Ssmj5b+Mc7uXOvODxT5Glssc0INXxPs2t7ah6/ylhMiY4jFv
S1V1TAjkycjnwogSFidIACXvdm3xsllBU4Vs3oVRF2F4c+YRWJEA74DURZNfNVYlAPnLktYpTTkD
1jyXKhf95kKYxIB9wspA5x2SvYt592W3cJoTbqnn/lN6cdlP2CaKVcHfVGxC2y3TJdplN1VBx8vg
is83Vs83zsxBKHS3UzCVAr8yZAmaUIqltjJ5lBm3cHmO7qRvWa3exZOydSHDQXeZJjCw3TIqLb61
29RKUac/paS/BN4M1MMk1VAdlWYWkUi74jAY3EAqIyNTApp/VlDuGfF+Wnex1Dc6UCMJkvP/1W4N
/dTy4bj4v+zXa8kk78NCPWFUQSIOvdgwmFfw2HvL3+E2+YU9IblauUtBA9ZYngATBQnROu8cKbLl
Q+6uUVRKEcDCnTneqzlAx+M/8LCIzR1jIg==
`protect end_protected
